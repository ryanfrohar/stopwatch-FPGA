`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PRBNg3KyY1TR8yWZsnJnzzW/dEsrSEDfE+1c6Hou7GiQUi2ny3LJr10cVebRXHTs9QGvYYRTSSn8
Gyz5sNLHnA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jp7GnVDs4XPGehBIKJsokm3xWBjOSlzqHCc4XQDu66HQLxD0ZCDJtK/0K8Il8OrKOoC65joOn1l3
Jor/QFU/jgbh9u8Cb2WE++syJa27o9YGvAlnaQpkj+0+N0NSqwnZUTbmC2/vBRF90ejN3z0SxSuf
7ogM20Bk3ecQGlrM6Fk=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
C6JMRfgIV+Sc/HUYaNdQ7GIkz8COMQi8XUszLwYumZyMji0WWhDsAmhdfX5HH8cQ2yEACYyrTdP/
TPkP6isgOtKu5yx2FXkdBxlX4T/RYb8TFzYCouDdbbojP0Ri3EnQY6Os7fU6/Kh0RGbHNIurolFP
ynqKAqHwVx1foWG/fGE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Bfx6ABSTmJJG+apj7DJxhWrxKS3DSF5eBFzSfEJkgmzGC4adPP0+EtlS/8cA3WS05a9ZnMSU//dD
6Xa665Pgb6piwHZmJXNDVJXTPEU3BZXO0hD4lShd7QESdtDBIjPVNllsAMr5ICT9aeAuRZ4712CL
OsJBlMyyKq44NbiGgoZsrvYB3AOby14WleukeyrHVRqOVOJbPwg9fW0vsTdksfdW/S6AUHeuZNZw
FQzUlxYpG1/ulxKJRSWGF2rVs8INdMkWKU0mQNfz8Fbu9kCy5+qtyDgko+t+9b0QOndyALYwiMoX
plKql5/d/127rmaQfARfQyiN2GF83TwGN+q8SA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uN7qo9Y7BtnOroN3nCx9a5nDr+AspFVYFgtL9vAD/836ZRiS2NZlcBzHW7l/qr+zJHZIwdEJdB4g
XTacuGx6jN9qRGwxsjd3FKG3v3ezqTrcg3ShQaxbt4rb1UWdD0rGM6JHU9UjV1v4FGjdDtrez7nV
yf8TbYVAIjeVuwTKz5QV7v+K5d3durINdZF1N3Te+ED6whBD4ikRKDsUQ1uT+omn+AEaJruouIng
kBII4smDkPDmW5SZwbcgCZanAN4z/r3pZdBTsYLi1WIMAt49n8T0NBr5BQX7Pwecdwn5uJ1uQo5u
PtrPHwF/NzhF6ki63bIUN1am+XxZ5abQxhzT+w==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fxhZ+v8RjZpp04TYOWBrq4+/hxS3PdHwNldw733sowphaSpIOkexyA/fRFpFYgYAcOEJQVdGxlwj
L4vfVCeW2SSHwtR7VGPSbEIqenEpmN/BMJKkAqphU3QYmDdQQXwymCL5qvIaORVfIz1XLVnp5y+3
MOyNHjSIDozEwPBkzIs1+o3qqXij8+OqX3X3AFlhB2Ase2TBfPeBFWKpS/1dOAq1BfuotrmuCum6
+UTctjS5n2x+OZZxOe4vA73VwVVKsh8ptEGksrnhLVJ9Qp2EfA7FXAksUYeGRo3dHvFOeIvvledQ
eavcoTOBjEwcPZkek4i2nhhzqQQJ/0ZEfxZcnQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99168)
`protect data_block
t1qCZNMS4sXqf3n+c9+JVxJ4ARD5DE3zoKDNJ3U6q3EGUq1CDQDoLWOHaGWILWVLxrjF4H2C97aW
tyKLh6hwR6zw3GCg1D0/sMKUhZvwWulGH8W/w32Q3x9Zuv3PD3BfAcovBbypsmuYYgBYlELvhgT9
llL+CkWD2F6zoRu616RwE78pqMh4R3nEtI59pVeF5rEGPIXd0sy7GrXs20jcq+HMUqLR/Xzb2NzF
cIkjR7MldoKEuksVlaU7UXl8LrLj5KuC9vmVzwhwzLioJJQjDjIMjaYmTCjUtGNu36WSnbfWXO9N
Ot2Kif+5qLyoHMDBZ3THUArf/wv3yNWx+YpOjdEx+MUvC3r24qhIGAAOkdjZRD1tsIuzxyGAtwEu
t3dcixEZhuWaAZWHlpVLY7l20AjtYzHxAcEEYKRkc7ki6frT7rpeOIFPKq+26tYoKVvyA6bBs0pW
Ec0r6mr5xex+PeMIF8il/1zmcnak8ai5948JRg/og2ppSIRcjvNFkTWUtrUJzWu+DY8MIoEFr1VW
Dr0bSnYAtlQr9JAcXsz6Q8wT091LrICzKIgTgzdjEotcO0H0R9ZU+m/e+Sy0z+qyRHcOwcf8lSg0
KTTsUG/EIKIH1BIDFgJ9rDoeXpox644+3hY6gQp4/gXudVG24b5ZSZzf2Lsf/jgpHabhZ4KaLNA+
UPMqUCK/JLiuIjvbquq1TBCJKoiey9dYg272LEP9UDTL5DVLyr4RvMfEfQez9qqSTKya/3aQxfK2
S27eKU7dEd/osZAe2+qhDK5l7htRLkd/0N+b3gERz9LEBDZGGASzmwWuh9tIDMFc08r0FMVgUIQ8
CeEw0PYuZ5Ev+pRo0a9KotsamJ3+QIfD28LYavqZjPTSGNF8dMTdn67pH26CbY7wZrBdCGYqyOq6
gNBaIlkabUcW2p6l/JdUcm44l3Rb3WDd6hBDg/n4sKpzb7EgaHPa4jaKXOHtVBlA6sbG6XNOppv3
QJG0rN5A7+K+GnNB7pXmhQiqIhVEhqN2VQDiHRj5h2ZXivvonZFoQv0T1DcyZA1fuuDWSChdgWZW
773ZZiAzJt9dT4SwSnXSR90E81okrnh1JTEefVhdVIUr6OyZgl3VwbvrNXtDcKt24VkussdZIt2m
4Xbxj4kTUbzgqZcyVI/LP3Ob91MspMLjO+pL4WrxtxJhBvNuJWP0DLcl43Hh/3Ku30ROIaDEpkLL
N5YJ22+73ET1nLPJ9Jm3uEqql7CVcjnuLyRXUdzVhW302y3YlFXu3bm475A7E54PRlOOSpRu964Z
h0jr3r2nJhPne7jdCFB6K7AfjjFLIRa5Sf9hCxEUvFSUWHnWHA0yJAiQFnDLjUj/iVfWzlL9sRSA
lw+axcGfihuyp3qDJD7taxvhtoTrXUvUyX/asSP/ULS5a/xHA9JMmZbF8PmCf6MHzU59gaaeSpQ1
60TMm+JGjihN75nDvjZymZjLSFQEdjf+EhuScuGBdIquc2Q8eIJMO8aptEe2TL3TTWeDnKH+NLqG
N2dUS+gHH74Um3lGk3ZjbRt4aolQDWzc5wFHpgNrZjytOrpV/aF2EDdrWyjQLwKRoStDn/1N4JgH
EAHppxdSY8worJjZli28G7/qBqZ5Q5Ir0oU1z0qLV0ji0kPF1HN4ceNSsE9hQDU936DCt+kF6eGN
0lm7SU3SuCJ7eFAOkxxepj1WZ3jUDKbYc/AtGJfNYlmI+xpwB0mFKNW7KACzeQYgCFaWCiqqgQOb
vIozFuZpp8r8bsdoxphl9FJ9z5m6kCefbOXuEuGfMCiVQp/pjqzcZhFYfVKXERU4+JpZz5CqROdw
vkJqPI9AiKe7Mp8rGNyXZqa89EXVgClar7leNYnFW0FcGvcHEGMExBCu6OwIcTRrJGKgsTHQsPSv
nyb4H9kUqBbBdhZwGTXU64kBgEIYcRyOnh/GwSzQ3cczA3Y+ZpJw0l/Bn5LwIMFxPVEXKy0XfoGL
VhSk+h0peFJwTvpO7Vf6xZF7s7BWs18v1UzpeNcPqRcAOepmIzOyXRD24K4z8K0gFNBtQvveEtfa
kPwXCTecKtpueVyAK+0Da5xdexeFrl2hBENy+5Zy9eoMaWf11G8AEy+HQMVkqnTQQegrBCooNkWz
bHK8SDS1hJUW9sU0DofsG4Tn2sXEfuwESfzM9qC3PUpFEMqyCzbS3uWZrYDBoSemqzEmIc6WagMb
Wo0pcVkfZQNelLkqvZrOFHVdKFRgeUn7/tLtGkXcl1BhuJ0LZP9Q2RlnPLhrOtZmlGR03v7io1lH
h6rmZrnVILzXY9oQLCiE1tPY9TqrOvlY7OYGFlykS7wFD17IkD1p2H4jAaoQxL74VxsLb4OOOo7x
Cn8Gq70LdyzR5syeA3PxQ7r7NQ3pXXBhXLKOLeazVsvAs4hivoHujahadxI45HTrab6a1du556mJ
NUOHSdEEOtY8cbHGwX0ZuqpXC3oCX7sQFh39ngsxENwmGj76yq4hWAmV8j46DnU0CHZb4fl3AKUC
eFG1RGEJa5OD2mMuarjsaL+rRi2GmStPDcvxc4dp/gWWAWqPp/hsIGn1Nf6jr9Fd/0zRXFw8YdBU
jmr8fqWTW2RFY/NMfBrW+4Q8yZIEqvXABOIrwQrP1S4bfvzK43Zj/+NPXi3RU88nZpJA4e/QV0T0
V5YTtPURnnzfs2F+zTKEhEZO7y7Uj4QTIgophGDrNsVLZ0QsO0P6BNALJNYgBaxXX5w1XCGIcnwh
GYUmRZbWpfSerUtTGlQsf9LQVohRx+F5Ze4IMDErlAIcv1kbNUTciIWcrRd4yQI2kOl2rcZKW/8v
o1ytSFAms+rlC5jA91bqhq/5O046/Iga+cbqgbpW3Fx1d3+gXmpjYDCCyQ6Vk24TsB2KQPyGxwbx
3vGKpw7/bX1xuGgtCUzgAdkapfXwQmhDRtIUHrF7mW59uZ7ZvBwEwq1pc5Xu1YEDE+I47IMktFUR
I7tnjiUdDCiVNQJtOt/eniry808UnJbcZ1XV/eHUrh9XjFpaZFPFkD5M/GV6MW+O+afcoVQD7UZf
5iX7QzpB5k5VIJK3deIc6XYCWUAlQIsn6acRU+oogUyJpKAxY2PwTRwKmBb7Hjc8ykLwxYSa0Mmb
smFInTZQYTMIX7AY5Wg14c9F7i+Q2le3EMxhHZg8oZ2y3/RUZ5LjS5YFOVHOicqFOiK/yWBzap4l
6momphcwystR1rvnJ5j4jM4D+3utjDp2ag6vwDAQxEBqEqORGBwokrxRY8MTYybi3N8bnrcaDJXJ
i+sdLDKUWMH/MKEqUT/WQAdpOqo1mieEpAlqz09E+p59d+K2LVPvml5Ed3UIorvARfOA+a7kQlaA
/IguW3JfNT/1G47hOIG7kbGgnyA/ZAzRnnMs9ERyXHIJtEhFp/SuNqehRQ39tK5166PulGjkLCIA
fAOhNxFaEHHclLRGKjQ2BSlMhpvTYspjd4kW2s5bmsCIjYvlLrnp9UNkYHfe9vy4lMgf2A7csBgs
AzYktGscsSKsDRX4ZYsfveOVrwg4txdT8zXLHndg85iXnLTXuWkvLqu1nY3fGpHwusluE2QSPcra
FltPlCPLJKnnOjxYIiUFMvHd+QJeKwuvbAJ9N90yC1uNvnwDJyRJDND33AT8I5f6ygD1gBRLS7Hj
6ELLk0GCrHTkEvYbZZIkDgT7KRGqcPG4I3rIzUDeNtPyciosjhzR+QhCuOu39sD//UDqjBPH0GUH
VTy64Jz4AfkgsnI+lVH2OHUZvtfF+sYDRd0TaN6R9wL1oNwtYVcBeESyys6ILPDqpU0rtQl5Vpft
GtDndmkEOytEv8TWnmiqLgt2Lpj0ojj3kh9RLIDufGE+Ye0E0RAEwrV73daRdWQxbcNLAwdXAq0K
wpVWxLKR4lomgk3vcSKSawYa5hY+RiW5gDBkgygnmhB1pxmL3rtYXdd7y+Vtzv1E7ovOm6kSKePA
S/GQ+labiCUgj7tDts6Kk2/fC6LiyL8UCrNkCxcR18Yw69xHudqm320F625Tctvk6gsVc1Gn3/r+
brRG+KTISCB7nzevt71nsRDv9eJCN3rE/aazIRZx+gebh78QQezlCkMPQJXJg4dpeFDHDmsq5mqM
09KT1P+QxnxvQ8lOxT4z4eLxM2wCoGh2cy9r53pfnf5Ayt8GePCyy8lB8Zqn29YhmApfsDuP3hCA
ltABXpMDJZjlHq9X7eh+8KqCoqlwoQHV7StNJcE7uxK5BxlLvevOQaruMP6TcStumqUf20CAElBz
6JO4EMvQpWDa9LR8SZp8l2aMJWXkzg9diLB6xTXVOmSF+GVsvjP4d8ArnQxipFPyDTNkUYX1Kin9
/PjMxkp5z9BJdiFNlWdTH7rHsYvxoH4ZmJPR2f6HkpmqEf1OOAdVZdf6LN8DVP16ZWRzTmco7+2r
iORRm8f7omgdYZO3eIMJTsSUpCvO9ep6XDiciJ3MDvkFgdUvtbmKAOqWQgF3f+AGgc9KwlvCSs2t
nirIevD7OA7dJ3JcdFwdPMhbOwabd4ZT3EZmw1OJ7FPP0MtdUBmU7R0KmUpilB1qGnAgBbusRU7s
X4skU8AMzv84KZVqJlk7YNX9C5O4gywP38NkVnipCHophOfOF7Swqb+1wj0oEdkYpXqfXvEcwAgJ
Dv+RGVA1C+46+x9E9NLtslV2m0ffXPZ1f9JLD1EkOC6n2AyePcv26TW7ewyF94JR9hQjYSfwygFS
KtVWiJnrdgdF403XxIqJoKX8CzVcuTYC6trwAB9rtM2Jv5ybO3IgGFa2oDUpHUR1FPSACiwXV9wC
aqV+qLgmXXuNsqXaewEiFwUNbXpZQ9K5I9FpsqKuRg3VKxqXdeKNwpZLZwOJM9/V27Lu/0cCGHmv
sz+aoA8KOBqJ5qbkAYmsoyoKEocQukrW1Nib+cmbl/RofXfnmjkQV6bj1+tMHkfSUvvYiklobSaC
oOIa13j4GOpNIi5SNR4JNiexIUKLg1Y/KOsLcFumcnd1Y1zxlBUE9X1rV8asoGFnhYd4+6IXzzYI
XF+qWGw+0r+AXI0aKzGFi+qe4AyLMmSXXNos5Zc63pPtO2VJToaOH7a7IMrLUFIgFFgc51iIq/Ll
5axkc/pLigX+4v3V/Wp2DwmJ7PdLOPwTH2xHq0SDBsZQLKIKwdYRTH8I2Owzh8DiioXpTkljsIOA
O8RZSdkDiAvWvB31bo7dK5b0j0tKO5BboNUfu9BsiBR7qMdU/TZo0QFVYckgL2emUWJZbCtZtrPx
dvw7wsUsASwMnlgONB3X7UrLCNDJbuW5Nm39wz5PVJgeZOiqWRUBl5vmU6qY2JA52BamZgTmeqF1
IY8M97ThERy5Xw8Biwj6hHfiGPM6BO8tVOVY5cpz9ND/X/sbxI1T1U+HYz639dDPgoanMmPOZadl
zc1vS5IAnXHei9QTEEM2gZNibR78gAGPQ9D2A6uYM7WKkYvyTWuOtgkvA+AbFa/z3LtISRe+UHzn
cZr+BSsd7c4P/PFAQYK6fC4MNp58ilsaEgVE8ki2Vr6zqARaSKu50A9dVJUbGWDEN+TLzLRJtPyw
nlyGbQRz+z2pB5nmmSxvCG6jwhLBZDlE6xMMKEkbxSgIbQk8/wm6jDnK1sZ/W2guxwSrEPTrbEcb
kEcTa1rm1yf+9y4oIIUPCO7TQDjzMARa4R7JtfMohS/qdVmsJYqu2BbpuMhDq+GVJnn9ECUeAhAD
N4crTya6oMfug3fzic6q25v4hQ9dUs6RlrMoZQiTQHa/DsrxcYG4sdwLBUL+mzCBVtKYO6pWVhBL
3ngyFdMqhVKRYidq86JGqZZnOxpWSc1OKGmUwDwkHgL8i+TGFt36PSTD9Q20IKFa7pwqU3saSbjh
FEJhsQ496bAG9EtbUMKpNY+V5Ivqte4YEcCkYqjQK3Ju1Vift47xPjFXoSlppVh197oSMsUGXCR6
mhsHIKHXZwqhR+zNIPHqXaax01MOhlMis1xJkUdo6wLGZFE3T/nke4tj1ez6id+UcsNHKoNkEp2j
nWdLR93CuwYyaDgnis1kkx1XAq48w74DEHR2z5unfBPZC6lfrzml6yq1sH6r1IWO4RbRzi2KGC9O
5rKXsdO4XA4n94tFTdqMAh1uxrBVFwNIZaMyRkjDqHdF3TPN1nCjTnrJnGSqKJn2BDyx8IutPY+N
UQGpUQgnkI2F4DqeQ0JupQk7n4Fy9SxcyfG8B+mmcAzVKXrZlf5EmAJT+i2v4SAqs5TT7n2eIWPp
7wcJtNOb4vCGyoTexbnn6WFyKkKc+EvivmkIq+lhm283wHlUJJN5JxbfTVMur+9S0WWloZYmAdhb
fO5L2X6umkevlZU3+Um9Gce7nlCUuUmEsTTLCWYY+EQnZnymLkh9EvLjKBqjxxdBLfapRQg7ndz3
dHLV8JSNd+HMPDWvUXNETIDIQ4mTcgFgoi5UnW3iSC9JRgfYwKzj3SSBGgmOtIYqBoTckhO942AJ
YxNu+vI0LWh4NIw2Tq7waYUNJBNicyxs2KlBdx3cHeofNQZjFRtHsWNzfvmwW2txohQwpxk1lI0x
iS1hYZTc6OZqagGDq2F6CocmOFDE2E+9FCuA5zb3rWu1O20loaufSj2GIwWfwMxV+WzbOokFOQ39
9XVi58XYMb/1nHzZomtNh9Dr6/7w9nTASooUEDm0dlj1HtJ6yBr4YraFePaM204OWfxMtK44NiVs
Pe4QGqqZ9H6eguLTrzN9tngEZVW70T6MtXHbCMGs5jIHGKBdsBgv9mgtWw5ciYWmfiyUgMmJ43MN
ruq1ZIkXAl9zLIt5BavHod6EKZ7cfHB9BvbBo5vG2WRgmWtdaUh9ho8uOcbBA4JkHh5j9N8Ozr2y
uJDHlFIfat6gWemQCtriClnAhbwBPGJMnekvCSCmsseaxLcjfXuVK1OD2LwR9toh+anlXONRh3GA
HjusIhxWH7GujpI9qsHlUQK4KDs6F9RbYcnDcDECf5xreJDIs/Ok18DA1KPVcLjInuYCFy0S0J7Q
hsb3vqWRKcjENJQ1vJWS1fFwP8fRPuKvkpHkODBebBOpwLofN3y8y5NTnL6rcsVcKE7VZ443CPA6
utKQaWoqguBpR1OJbuboYtoQ9D+MWraJydiCA9yHHHkmNvyz3H3RMmYq29JWHxEYW9ol0AgbPCSQ
IxpXgo9cbDIRyDMobE5yAojXEPscZybzBD0TcQTYPx1rWivEuRLDQ9NZl6o9h5ylf/tmqIToKBle
LK08RWIJ22XlQRqt35bTRz84y/2QMIXmrytbzPD8kHwu1RBfx4F2VdYNIa2keEjhSMf+7gRf8v4b
dm2KkwmT9A6SUoyJ1K5NmrlV+QdRFeCOsmJp+lL/ZHtFE24WBo9wWbArjLgbQ1zLjOR6pXk53yzj
wjxkrHXzpZQ4ZTMhF3WOiq2xuVyRCmS+rNkCf96av+jpIMS/+FnKlu5vn/WBXh2ozLSsp4TH3d6g
0HmBt+exNmj/50k5RjDw/q/v7nxohBxf5cLtYS47qklPybAi9XmcwcdeBsG9UwFl+y2IXRut/g4A
1Jb6WS8sngtNXGUiL7trqZl/fqtmmFblYzu+O1FycSDHIGP3Mj0vYqQVVVaeVJAtcoGbtiDxWAWo
x70vzSfMMpJDHuLkF/2YZ1wOr8GgG4VUE2JL+mCldQbnYBYBnhk/yPKWH0vZZEWpQrPWEejE0/q4
kMKVJyySnW5M6tifpaLKIqjMgu9/iddyi2k+FwGxlF9dB7hS0lhb9l9BwTco2bEV8tKt4bKS6txy
lHECGDm7L7sjwnziJYRFvS+MO0rgINmIryBO+r745UBo3Fgrt1JPYJTpK0yypRT1CZ3ZnnhlaZsA
SCJ/UjHwOTvdX1nr383lhwWoTRy1xKbCTiSPG504QBTuDM/i1WnfZNGtzfv97n88WJTcF6eBkmr/
Tq3J33snEiDfrBLWUFzhhhXQmx79qZ0jnflUmd0GCe+oRcNmdRfclQuWWj0VBeR+hHoKH3502tHN
aih6X6pA9pjowHKFhnX7FLLsBVUOu1/3P2D98o5aoau1hCzU56/JBV5fqbhHm/BZN9uc7kE20xBu
EJFV5Ny+nRZhyqzlA9kfgwu+y1yP9UE5OD9/APkpddEIxZDgE4yOHFO8Cn0EkECdVwP53ANq0182
VTEX6gVGMpWRmbVp0j0pZdM0eZVvgf5htByIgqZMbEiL/xMXF89yRsrAinQ5ZnO5cAI+rpFBx5+y
6Sddv31hBBZHiBPvXNL9eedz70eE2XpTYjiKVsSgCt3TY5zpWuzfz23bo3nECxgQMo/A9a1XOUB3
1b2B/O5539PZh6OueZSrfkFBo3Ph5oGQEl4hQNO7/F8rpZ62304laxbkBS86YzvwanMPw0jt6wUr
sMKU4P5iPNTdv/tk56K/wk2Im3iyxDJ1sx2Rgqu0Kf2NTBO6++8+V5MkWBCnjeuUENpq9XBdSqw1
VHr6no5IWu7JPN+77WuKpYLQnqVBQT76IDCi6tCHjdE4qPimb3yQChlJIkA//qpRvWQRW6ExAWV/
hTHtWgziCa2CDv0OyBUzRNPYXZFtFVK3/PVsd0CgvZHk78ob1YEUyFn2fuLp0SuvX+XQcKdLn6dH
tq9wd+rxJ7gaddxgzCjwjM18d3GBMV+15QpSh8VEO6KgEmP2py+QwaUMhe1F+2Q367/LZ29p1eiO
owC0/jyqh0UL7lgdD0o+0yTv5oreVgk30qi0E9lnt3nzbfqKo6T4Jf/tdikK4UR+CQV92MYYiQcq
RHoe4hBg4ZWrEyoGSjA21EtFh5C8DmwKjepyTFE/2y3a5HF8k59AJBa2BXCeRoS6qiY9KQge4Ckk
WdI6gXjUwHAH6LCss+bM/kXLWuzWTVyxImL7r9Xa4vpP19B3I5ClvmEpgj8I/KSXzNo/Ag2AkswY
r4Q3YIRd2yfXtOegYh58Q8zEsWtZvt+X9/vWnTi1RegsKkXED1a8hel+HGsVTyEJ9qe6bmTvnNJI
EVmLMhzPN3PFz5HO1QV0hg9M/ZP9d2maBhbNfLsIloYrtuzZq7v1Gj/eXd0I1MdXWOJMcIWNA10L
ufz4K1mIZktgXLxqGWZLOneaHrfwlLN6IYCOHmeyX1e6Fk8nuGNcyW5gWSiGaliUpC/fBhhWl2ZV
4Yx6jGNWmiETZ+u1rjhSJYU3E2X6IWqhzubSrr1rTdlBHhtpsW7pOUwl5DJeQn9Ng2bpVwv0cRK5
2s3up3z9mmHVAB78649aR0sWJufGfnU4EMc9oHy6huPcEVgs4F390fVPL0yiEPY+Pk42Gk8wxURk
y5P+6hecO7gtjsVcB9yvyFsEdPk/TVQYTp6qWXHu7h2Ow/LfJu/Cio/F/8MOjPtSzxJI43P5sYRt
fAXSM1ln3WW+L7TCUikO8nZ4bft0M/vPfP/BqTtjz7wQ7b5/F+8HWOLLFbhmCWU1pIu4Gf43E0zh
tw+1RnRKwqj9ATBC338GVetzK3u40g0bXnpGVc1leucM9jOI91UsVakrm2x9QQlsyV3sJiPaedOZ
J18a/I6NURlbZ9uEqAnCsEussi5UXZU4cM7ACeRDtGKxFU05pGl96WOVG4LnnofVFb634EaG4mJB
hWjMHioMkqDtHSFdn5qHIyf58iMCfEE601VbCKPQhhP6429dKBAFdYzrG9W2LvjeE5U2m4RPpFmn
KquM5D2RHU4+ZvHAKoi/O7Jvy7IdW2PNQ9FKThA7Cg63cb4qyWA/06pe1xct4Qkfnt/f+A5EmEFR
aJypGSa9WWPmMvxUVrzx6y5GRcBIbKzcbR3LyhJ7kbPv13MUZ0uwMtrCI44BFcigrIdXEQ5S4ycb
CGsTUmQB9HZiH8vrluwqvw9fd7waN1SU7/APA07yM/U0NV/NJ2ZkcqKBNyHfrf/FNaBPfHxZsVai
mFefVqDdc/3Emm3Jmu+9g9UVLA7pqfPUj4+tY9JVrWbuYTNe6wQObmILIWFM5HqLzcExWscfthEP
/Pa9j7LGo0sWaK14m3sCzknjGIhFpzdIwNlfHRwY7RLWDyNmHpbzUYGCk07lker75vzk6GvZ8K77
lXzN3HVagx63HXVKO8V67HTsnD5kKkc6b6Njb+bDGmN4zI56YQ+/kd2bBWydYTi1oOh1P65jvzJP
njmyQyN/HAl/bQ4Gt7ABpvf9yZd2gO2tAlOtJ010/mYVBLEeBJMGJxAR3nXgMgFi+wXkJszUPngh
5/yIVBylpEtB0lOLyB3v0aud05jhVRw6N1yY4qrjYv9GKkHMQkcLPBHEijqoFLYmoQFIALou3yZL
H2oR7C0wmMwXD5RwQsPkacD+kbGgdu7Q6o9VeGo+1ca1yDFp1GMbN38ZmBCAitzZiMv6UEXnjzX/
oMiOxK0aLy/gqLc35CMR1Zvi0DJHlAKGXdVDiKnNDDVNN2XZpYi5RoyHhLgTNUpQ3Etxvd2fn+Sg
93Vb+K0Wiqy5oWD38sWKfN/L0/SgQsPXexGS8GYxCdeRs81pIYIOMaaKmjtIlwcAtu9sKsKOhCYk
s3L/NGMTu+5smYLpQ5ss/CqTR//ymMDanadbTCioP3evRPdzU62UP/Kc7OZLyiqrLgGFZoYiaJ7w
NgcysR6bjItH1AYTgG3BQ4ibmkigwHPGpHmtPfbzntmyfw8Z8mVjYuHU6cQMGT/Pc7nCa0LPtvn3
7gYHTWcv3n0HyeOqVopO/5n1MIEUnyYFlLEmNtOzRtulMPyc7ZZCDYkJGylKUiPX4st3gSzZkMuW
XznnAQyrxTSKWKl2XXK3BDwwP7wvtmRBCbCaHV4u0kNezBU9kUnick+NwYE1P2KWWz4pBiRlCyme
LLj+ND/EdA/cELB7A8EfS0gVQSoNQgBLhM4mdogGQvkHFR33DE68VKeu08VLuiHszSPSX4tU5i58
TCOGr6icZkzRzVi9kjUr4ZxGfeFlZM9tOXz50jaQL64e7roeuS5n3CbX/2kywKbMiXWIbLsEZFQn
Cid6IZQoPo2E0jSZxN6hkh6GYdV6wsma+jHSrjDwuxhbUqldxqNRt6JNCJVkxnUhjz26l4uyAdD/
CuqK64HTYzM9olSP7RCoAvDGxmOt4urV7SJx6EFvL8dGbGhu1KvxQYiDCbpOlXlLR3g1d+BL2mOM
PadUT/W/i/pdh6ZCjHDJEEOYyt/HgVwHeQryOrWaWNcYmbBgEbtqdaxHxCdYczFJxdikAeyfchSI
Y4mWoRv5mAADmB7RMUOjUzE8btE96QXUM5gxJ7p/SISwnsSQskkTEiaOvw6SW9v7VujmGMO1giNO
Gdm7ZCVY87A6o/zxZd3G1+G89A8zVFP00oZtXZ4YbIRReRgrDFE9KbpbDpmj5/yYkN/JaN+d12lz
5bYueRKpNrm6EmkTLp96gUJC4QNsJguT75VF5DLwZ124U3B2gUfWSRPTmhgLvymrTWCdrkyuqRUR
oc95MUhUqW+qF6n+iJOnLWgdM6UjZKd/4/lSMJcq0lF3C99gdiUGsnW/12QUG2z4tt+16gT+EQs7
m3vtSupKNjPH3QSqY9knFHK1p1MwIhcONW7BbPGCdOtBbKKizzB0afpTEDYvAq0U4d/q0WtuRW0l
aHxCryEMhmdEC1z2zggMo4T3OScWtlUgo8yEYGnKOwy1i1mw+4Uc7Cq8GIrZOHjLSJY/ZR1DwFbA
qGNgQQ/3cqpDlzoF7DZQOegUefz9UlFfHuWNNRZRGieJ94p8Q5xq+z4OgBu4n0MEZBxHnZ3K+hua
PiiwxSDisFzV3uxS2fi0p/PIwhmpEDo88N3j5pYjwvx5iPbhdCjJcnmrxMGlG9SUPegulV2E1Wgw
Lav7bXkgdhFwPA1pP78VYecgidFPjHTpFaSjWhCljADuUx2UIkJoD3MljN2OabcwpvlhYm4Ofa9/
hIhkrNwZZ0MK8vOItvUWlFrYIoZO2NxHdVKXzbpmNtdg41Eg0kkKQI5KywLNOV9QiQqvH92QPgRQ
pDuHQlRIECDKhM+xhxcMYpbdTiS6IW+dLYRxqF0XjMP824J2WauRbXe+m/Zoo7KvqsBXGN9vp1ay
icpT+Ug+YqtGvmrdCC/cITovsLyE/3ARZ136XedFcY97rEvaeZV8+lFD8SJ5vxvqR/aYN5LqUrNl
sv8QrrQ1Z5kvqlN9srSZ/Yx27heYq1Xf3EBl/+cYoCCuiUNEj8WK75UPizR2I8mJvJcJOuISutvw
OMNM5bmY98xIznYSl6/46MdQ9kK/rES+AXG5fOFZrF0wmc6/ghDzmCE5pxSmUca7+Zjeu+Qt0I89
fYIa4GeCOkhmRZ8veWQM080/WMctp3DK4N9B80jMEW0gzwD3Glf4VEs/+7XUaQuYa3jsEHivQMHK
H5LIBCLInhMsuDT144wWRJrtMMa33HXwxnTwbzJ/sacfif3nZzngsb5rWK+cr45/w5TKMd8S4lmH
O5OT2qzJ9lrQhpWBhwn8YV5TAXlCm1psyUNY47VuCIWLDYbXtDhpQxXw6S4UpWAe445WsW3yuMG0
fiyys15dDacqb+ZvMzHfdU1vltJQaaLsPfmV7xr0uMjXTsB96vKghbrlSiS9Z2jF7rDe/5Bsp1YK
1OxjpboNAggdTDrraUqnt9U8gC9m7ZugU5+NTesD7TLRtcJlBa90MgO/hr7n3iEDNlM6JiHT+lFb
UFJVkIdwhBe657ZTAzhw0TW85Taej33T37OAfuzcY9ay8psUx1pRyTr9pBMt8QH+vprwQGa2anS+
cDhMMHNzTnjowCyRNCvt6nkJ6hS54K+vkS+oHHNXaHTbJtFdF4aEDzBA9okmFeZdnAXEKLZOCxyj
1haoGstaJxkhgJsXg0tlZF1OHWIUa+unk50cxjUuscaeu0mGTIwZqdRfATepQdRdQmIhiRzOk6Cq
OFoNLRg7dkSCvsYCL/DBXn/ikFSWXzIas9Oh/rSIbVoqm8b96XeiUFa3ATWLVSzhKGCitek2SWUn
5yNtll3dITOA7j6V0PAsYs5sZkJXMWoaTdrpvVa/ngh/cvtrOVOvlHlj266FIuRd8XLH19Qx7sMZ
+5ethGs6iwYNLlpkbU2C6vWqCu1eMC0bvU0k6oj9RWYguQKTBESV6+Y18gRywbwSTJYtBLxfCtSP
gM4OHg5AiscVn9qY2FtBM09kYx2SdlkkG6ay0RqEWNLVwxVAARSBOmAeo/6Cozb1J6eGs2lpJyh0
x6fahBWV9kj8llcgGoWgw2q5Uy7pEFfSzN9DWTw/oQMSu/NArP4c3Rimn0ra8cC1JctlIkPGIA/R
iwZ84I0L/MbVajkayWUQei/z6xofbxxqZJLfeyJwXyF9OANa/a9LfsexAj194Cr1gOMt7weUaehL
trkQoTysNc7A5PA/YBnn4i/TctoWmxoOnLvAWdNWoepO/QmLBgRcSc5qc3XZhfalPkUW6wJ8diyr
1jpdYT9yMP55cH6wQzVnoZ64cHeKiCJMeRM/MOR+1s2u7iJSYY8wFIrAZacvHxmk6h76fHKN48fl
Qz8ZwjI9NfDOk8ZhV4wmUfiJ/JBM7R2prhnthXOeazJll0NkflFWuUJinHyuK81nYjIQxEfsa9Yh
HAOP99LFCmNUYglRfXRECJVV3udIu7TpfTFHOzVvSHmG6apcmAnC3W3zwu5m5TqmwHBF3vXBdrbX
qvrPATZ0y/iRurfLkGE8+HWCE2bVEoHSpTSNM+UoH89oHhA9izUtvc4E8nH3O9r+3tPGTGFDQ+EZ
CMEO7H7k09n9ip+3ZKHnD/GXk4XJotEFyhAHbXsIll3ckUaFwJgHVOkGpliHg+FPPjVJ0QgTjR0O
DF8c7QUA/8qMDrPwcqENAkptGklWruBqPYvbqzUhebz1IBwi61fLHLAKGxC5ZJPmFGuTrasUG5Ji
/oYl/vOlAkF4rGYyBfr0Ik28NOSKUHyaNPoAVThcoY1uTJix9luF9iqqPh9m+C3mI6++BQ4ncPBP
FmL5oP3p5rCCkdkmZCwqTh7wdFevfBZTYJFhiGPfKcvskMcPjqaUaR8SOXiL3Tv7U1+pjMd46lZm
J2SBk59QXcLOVhotBA2ihTrHpmfRYNlKKP6yErB34jCXKIIwY+Xc7sMxgKepQzCTqnckpNNk+1o6
s6+WoQXJ+Ix6/U4lk1ucBFXlmFfpXT1VcA192cFmSjt5vqZ2MsfSi18BvWUQBkU0JkTucf7I0GUa
8QgR+cR2H8X7L3PTuY6B+BLDpyqjLPWSZrpCF0APLU2T691lUVsGJFDJd8rdE0csvNH9tBiYQZVx
Bkq7fYMPlyFEHFCVzjfrzLUj/VR31r76Krx6LVB4WExtT3uFzseqIuS5IB0tOEcE8ltZn3PvHoi6
9eqeOL5bgbqatGghc/hxzus/Xe6qYMJKj1TWtCn3GjfbIX889qo0TKg0Ls3cD9OBEZKtoXYJlYer
gVgNMJbJqp7HhPlCKVegzmXTiVvfMjbOq70/4jkCtHZ9ntQttVsmBCH43i2FJf2w/WtQ5hPc8mIG
b3REXltLadJZ4gvNQ8c3ZPhdrl0a+yn93tpITJ3L5MpeU/wwwwdsGDgbUzDgtJnrLLwKna8ObJgR
KcW51IHNzozQfkv7rMkWq1nmamkoiHQBTH46htt6HCIt22MVr8VQwZYstRPG1O48W1b01EmY1cjN
om3yRZpVQFg595bHGkZiJx0R9EodHuXRdmfldcqykBHjkI/Yjoc5iUIWEWA95jPVJkBLPQqH4gOm
EwHjU4U4Mep8VrixMDXwQT6zXm+tfy/Uw/9eSI3DIln9yL3fY34Z6QqnuQlkc2uLVu1fLQkd4i94
+9TVEudKxEZXvmggz8vA1F+j90Ywk9uw6OstfWkfiI7DjzPfwp/UsgvXAjBk9czm1op0SuGCLvz4
JOJaAJ/fGw0Mt5wrw2GlQwMwBL/E+W8ZTsxofyihXrtryRgj9u5UPPNYlP5Ye0bmrffevj2/+031
p1BKvS6YOYCHi8me8VUG2b+/KuKCHAvTn8XFO6yd1QRuravqafUA0Jqi2UkW6IKXauMXr/rgAvdV
hbMprZXrUpqjRy7lEVVNJeDH5SIqP+deLNebk4znxguGM76Z2IxHpZ9V+BcBDWuGnJBsS0aNQ7wD
l4pgheY9FTo6rlKRYIv4+42nBVi068eAUjJKBOpeN1B28AbOu68twmNvQkc1clC6JN/Z+xB0FzuE
Q0LhDdqzl7LgCQ60QZ5CFwX4xHWl8o8VkNGl9JtQ/nXH3n9sVV20rkS/jA1uNOqq9kqps6YDQLEe
Ob/MyYiLVaUjthVBaUdJMHjLhFm+SslhcQYNFWq0Aq1rjLcMqi3Zh+vSgmGtlfkiW22kFksMGS7r
8lKL1W8T2gPzGQ4veKLlMntZGqlPRoK0iqtNNpJk8D2fmvvbjJlvOZICojbHJsjrkccSRrEkDIV+
znwQsNZpBm1IOcVlHA3HwKQB0bznDWaOTHrsgQWkNBi9+ZjKn6VsUbTqHBunGr+2vGAjbH5RBf1f
F0ciCxw5jWevWeIShNjYtdwYtgV5AUd3976//7gqDiaADw69nVlveWdC/AE9oz2iLBHnLwXWkh9W
sgAKIQGN/wD/xQ1VfemdovoO2s2M7AH765eWdMDIHSFZNbdvUCa11VtjSieu2atShgDCuoJeA6QI
+aDDLpR//uRYt52qRF8uyVIlT4Dp2kglIJCodR7TfnmDcI1BU1k9GlN+nmidx3ZBLOQLreDkIdSh
5ncUmgjbPOTUg698YgMbdJ1ZHdzb80OOr2A3qwW0tCGWmsNJC+bAqADYOS0Nou8f8TzWuVAn+NWH
BAy5woTgYfQ5uYSdpfMY+kyzX+S7PO7V8VbSfUo2uLPaZ0b3IJhGqeaa3RR2/z0Wn2AqHrOofAAJ
z/ayn2T34BWCyBCi4cI4hfdmez0ayMXzhS8UTmA507Co1t7GMhJXTTGjjpuORRYATLl0mWqkWrjV
WTjqpQJz6e2/p53VP5elK4pQIePgdw0cViZmf/yxx1blAZL5a5nqivbZ5NeSjwuVgFMvQDuJPAUo
Fh/dmxaucFJFqNt1a9ydTsc8AygHaYDKPZs9ZqIJqJdynsMN4yrse+EkWlPw6z9Jao+NZ9e/tkwN
3L9kMovMlCUY1VQJ8vEJZPkIByQoqvsq+k8sqDD/QA/PvPh0QGgZfik0pfYPazZCnGKekRGGhWu6
I1Ei9cXpIy0DxPV2zOn6c0Ry7vSBNF5Ngj8CJ3RlsMIbQPx81MXkHnFqsFl70uvJ0vxxAIqp5eA3
+m3GEnGQCUuDgTNaY2fZr1sF+HFe5mOfvjLrwWQ4WR7nc/Yoru8S+N7Ehgy0KuDwGu/hyckEHYzQ
hnqWIK+65m3+DgjbpC9S+a+sVBHc0LUEPsAwzLqLZjPtPGP10VugfTlNZwihGwPPBR+HSoPqxW9X
tWqAyYYcz59Q2BuHYGsvQF9vvvyic5kbQBJJ7wEJctsZqR4En6eeGjfcKw8Wemji1hxbo+AXJszh
VaR4FFsYAsh822nND47lC36iYJ6J7LquCCwBP/ecLV0vgLoJkS8t2wm+gyOYUZs1M5En1y50ODQe
3s/hN2+0vndsGa7HxOSRpLRkshR73oaOToR9ghHq7Vxapa7ojAdXZhFea8kLs+7l920rVlPf+FZa
0RPDPgDPnthZS4vY4iB4LuhKWzDwdZQkiMo1gIM8yLP556qQAzX5iVBzt0ydTVMKLipnCVeOJByx
IDuuTAp3N/mhHwZD2ONksECd2D468RxA7zWMSLTo6F8RgK6LoRI4XjUlKFMN+TB65hnywuZcn3rG
yPsxgxK2JWp1sWvmi2gROiguCcHV/bRYJCGu6kGOKub1+0YSzD61mblITQdY7P90bbUOuYZMvapL
iOLYOHwTjUSd1rwWR/wDadqI2zGG56sj7Ide+DC1OzClsU+oY8c4msSWVGYsHzHjcx5YZA4dJAnx
uAoiaKFAiXjVIwrsd+CuUo+Ee7vGcKD/LasLrPRHpIAohobDZN1OZqy6rWoETMwG1ZtarJKB7zUn
XAOWhfmvpvcsCu9oL16FgU7YyW8JJeR8ommAots1ycBPKNE3O6sAAUIXxzyBQPgK+OhMcrUFT6Vj
EupY3LehQbWaBYhusMmKgTA78HziNjKDYFejWxy89tE+qwSnnKyjBu84JuTlhyFnPrkfI21xzEaY
xqd+/1b+ypWgyMG81cRfGHpAhr6wd6zghCBsdXP9DjQ2Kn+AHXePN3133Uq9ZobP3mMmV8/cfGKA
G6JSy8C+00FbQpMVvA2ixUiMpG9BTJjg1IopbhFjRobaLu4kg21aOIxQBQDCLKzMsQm26Dg7ufnM
sZm73AST3uKh1LkdzZKaj+TbTtyoR1csHt3hSYYLNf+s3xLydmkMvVHqCr5ly0sMOZbIhfGbg54n
XMGH6zx5zKbFgpj7nacxKJ7JqJtoiWjV12j9ubReLDBzb8LzvK5Vnz2cA3nymleOCWOSKDNGFRIT
yrVwq4svG8Or6SW6FBgphXmvk9DBeshALBVygij7MoKpiwDUIKQKjgeEyBhRjpyeMDfJ/o6jOv9s
OaveoNSEt3qTG5Ic5q/0/vccBxihM4m173hoFUTh0s8IHVRbZ7CAp3qenDqSEZLosPfzfoMHdv/0
Y/xRmkOC+d/g4lWuq+09/9HEQn1SAY+/eAyAmJ5m4R9xIG+86q4siq2N2CWlRiFlGyGVo2+W0mFw
jH272Wpf0cU/d+pOtFyu8Xooy6gp/KjRbzdJpQbnA+bujaZ7gJ0B9HNyPq9MWt2yR0VeyIYdKD2t
aDTwYQkmGvgBQvzDJ0fD/DFZUHoKNLG1t+8NYqAluOKKLnooKOifXlczWepdo0+UoTKmIZ9GMOG+
405z9xDvYEXw//SvDcR2HqXf4mOzq1jajg25I4gsrEufAFhc5G2kX5AoCGXLQiQgj2wO27Kq1WQB
3ollcDV67T+Js7qFjR1CJ9th63YuvdRC2qE4S2wZnJU0dUAt7UnwRWa4Izby3UjP2Uz/uUJm4XZ3
O4B/WRwrTy5og3qpiDUWRsmktT/tmkD42G+6wHRyxPa1qinRW9IgqZDR/9LpCrwt9VAp3zqKtuEJ
gdXKPCrh+yvRP6UnuL4Fr3MkcCkN1iPVRY4fS6NetMqiKBB/PZxdwJzFnHSX0fJpPTZXNqOxDtIg
hG00XjW0oo3ZgwKctpSZXUqsAbMMR4gD5DnGhfZR4R4yCQ6TdcSqh5aQGMfc3k/q59Si7/Iadglz
bVwiCidHAHEf9BUoTjnV5QQbmxCEYtpdMup96Jz41FzyE8xMKxYeGGPfyYM3oWbWc0S2xdBDkBnu
/zqYhIo2hEdU8hqCESIhrQ0qH25CK8uLQmOrsua+ny//zDrzurRcsq0MbA5H52AsLjRaolEd5Tzj
hLtlz5sZAyxrClOchz19yd/NMqFSiWxdvorOO91oCbaMcA5IwagwKqHgGxyCxPrSlnfR54wwEoSC
2Rp2KBcaDIL+Us73wA/mYtpCGbcndq1CXyyjQQAhtBFRWMKyhmFbInG0u6mxl3dRq03EKd9nyDwW
lEHjwTj43VJe+xbj9jYyhu7Af1aZppAL3JFh/p0nA567OOB3pY2I4GdDheWqtmvU+iUvGbepVR+H
uBRiXpKQYtTgCdW8mab9aWBcJHkhD1nHzVvrD+a3pdXdu88pCk961+uAWLN77NTLWQgQ1oJ30HoH
EafpjkoDkvo2lo6CQ+S8e/wa9Pp0mW0EgLOlNJwkuUPesejjUfBrEJpRBPpIY8zSzB/RVJ5Vgh1+
McGdZgwnNRWIjmlkX2tChlKGeySgg+Yyl1RSb4D78ZHInwZteSmX6PdplyaiwW3IMKYfYj7gOM9X
zk0rzitZE93EFfV5Yc/9ECUcM6CSHVmMl6vVIhTEHjjYtFG+Cdm668uCrCLtjF57o1MyYUR+A4lq
Ju/gFZbl0fHKS3Tyk+zAS0ww/rhXqNySwHnJn1pJWmJoBbAllc9LGqLCIPt/8/UFbse1DLBAdY3S
UXz/EKeEKe9B22tMFVBxgMZ890a3todGI0pKNH6L0LqoN3uZ+lJztOtFMRmm+Cs0EpmZF4IItSkd
ptYi7Kw2M5JDpWcvPHf1Rm25bzb4m8adFNxecUvg3PaE5Ahfwvvxjny7J5mjXwPL5OhATKWn7vPi
wFRTQt4/TdrjUZZXqdiV7OUFsjVVoMOlsCFNOxcxwUUy0EwTt4zpELWT2uVv2q810DJosM/s8m3T
ONMzhOjukZ20aj0UiTXZALgCxc8aSF6zEZ+5sQT8zauFdO75xuP6rUBHfjkN/v/xpPL54T2NTUvn
ca63+Rx6dumzv5v5tekO0JoU+jwWjX2b6hVVDz+FvPh+G2ck01b7MjnlArW04ivZLsaYTc2xrfSA
4PAeWOVM4vWuo9lxVuZx30dfGllihho0ioUWoEpzp34/XfyqQyLfJES2lB+Y7B6f9k43fT9XNTuH
71DLuMpepV+NZjAkpqBTXlOqgCEOwxsgFYlQM7kax0ry6lExJu5bZ+iNwTfU5Lt6fLrig5t5xA3G
oY9QORULw2b7DNUyVL6q38pMhFzGTEBEFuhGDmUtG7lgD1HFntaJydUx4wFz0UR1Xpm5Fu4GRKCF
FeMCvYNc+K6aiqSAL3mpPnIamXiwNkiq1mCeJ4bTjmh5HoImV4u/gwEDFd1dDDRlfqf/pZlRAEG+
/2Oku1l3K59mo7BF+fXA4VZr2NioZw9X6rYNydVdum7qfCGfsJDyALYXLvCHdoXbj+kCAhkug1nk
hcPNItU49PAGD/zv/tKMUHPRrqoTygVZIUMgZYBzo2W7ojigd+LrENtwF1yn8HGc8K9V9YBQtl9V
YXEJBeL2xF95RodoALkRMkp+UQCJle+dCEErpAPK//Cwhr7517QVOJfiTq+cEiCwF6mM4rMcOV07
FMgjp1EXalxNMmqXSE2ZZ4dZglUjolZpdoXlJtnwnzHmXP/zmENGJl+soU276WmziKPXd1CM4k4u
F3jCAal5pN4EnrOzJMbly8Y5lCBnz2clBFTAfdZXHw8dqTb37oX4TzycB/vIkrfr019e4LnxSKeT
J+weR71TTRoiFzRPWO3a/EoNrYQ8SqQBayBNnUBnymxGvWBe9Ekm/KNvMnoWGaLZmPAGPBPkPIUs
YeefKO+IFAeMFZmzo33NDmA/JvNiwUaqe+T2q08Wyk+0labZkutm0MsDdmX6dFcSPsHN6ySQphZI
n39fdSldbPSqk6iRp3M82L1d/kCIORGatPvo+0o4Jgp65nxd29nD+eqaHjV4ahfSDudrhDxTTDaL
Jzq96X1535ol7CXoyQtpSqz74BDkM7ga9A7UwN3Df6DiDzjpgglL2LvCTh3f7B1htA5nGELMZUPh
Fs1Q99iJAzRRQ4Vl2isohMBpspy/DhEq18W+zUlgnutwpe1RcxL5f/ccNJ/mJTogs52SRvL2/Sr+
uxtcatS1pf26zFVLp5ZmjQ6p5adNmHQCqYE6l1HLtcjEh1dbEsHv43yEbgBH2e1BUb3oro3LksD4
5K7EjKemaTVngEFAmz1CWRmhTVy5JIIcDo/Yb2B6kHEtRi3kZpvu7rCqxlbckfqBZTC/ywuJGB00
OuBR0hI1ri7u4SxQohnxx8dizHapwKPlnDApDenMqQNsZmE+LbvB+cngU/GKeNyAzPSBNaNzPKz/
CIeC/DoXspTd/foDYCVrxsW86LBZD80vW8F/mIofKkBTZyzdSSSLGq8I+MNVOKgNK0h+exTIUbhy
Jv+3iYpPYvn6BwjQfRy3tYSjwGl3mIgiJmYLQ+5EmnF9lzHbiGFYSmcZt+V5UpkdFpjnvTA2kJQM
2UyDht9UvFNLMU8YtcBHiMoCRsjRQHKXnNWixE+WPJlRlc2p7aWVmvTS+QsjroKT1XWMVeClT8u6
9PEGrkaAxfEutr1lL3Ht48Bg41W8EFjbHDnVW6AtpQx2ev8+XOLGlh3PjGwIgfNC1PGtGrXLDWty
dM426xh7/US1Pb3+25A+OeIdck7WAT1Z5XWXdUmKiqe7mIFaWNIPRs9gXZ9DJ8f0Z0nFGHBI3ot0
s9MDGyR0HZfT7QwC9+lSPjKelsuFaQAY6swnHYUOoEWTW9NLLUu4a2zexcJmcUG4vZGa8YgWD7Cq
+FXuxvpOgY/pzIMDFPQHBGz0XEhRxk9h3eaNWer4o3e+yC8hsWT53f7N3DJxY2lMQ+zzCZoaoX3f
X+mTqXg2TOvtiePEUxKO8MzljsUg2VQDemN3QhUBPeCI8lXP3jAHi/FcozMR86zXNxl6fIokzu8l
m6mjlfmfI4CpPTN9xhMQgNrlSYGsX9PA5aIfnUSGk0YbBKCTVIG9i0LGg/n+54swepifebjUTlV6
n1XacbtZ9PLEDVPACNLw4dioauF3FUJ8emErr+t77Jv0Lh89PgcnCSGRrAwvbdizN/eI86aAA1PW
WJdBj5kdOkZ30qjBxN/lRSir3niPu760u/MnttcweIdunUAEjmR4dArqYxC86sFhZ0sR2JY5JPz5
kvNx/Jr2XDuXZzTGU/6Fx1Vj0NuLOs+58Q5EnQRG0+5e8Zr5aiaYZX30mj9BWH57sDG9E4b8EqmI
Vq3HipPzizP9jToosRRA0ACKZPDN4aFKatRRVR15o1FeTReLxEKBFG/9wpU+I9HK+6rWvEGqpOOn
C3Zt+A6JQRro8Cg3TFxIKT2OIcB6Uj8JQbDVEsbnw7n8iyBdZaNfo3+4r4jtM/nwxMk5ghB0Ajnl
YoWAo1Xls4mNRU4tr47MM9RWAGLc9Q2kQCUGLJASZQ2Zu28h9PzBd28uaJUMZm0PJ9ri41g/jPt8
gFl7IPZbaWlvXgj8r1EQ0unpCTC4f2exQfyIKH6rxwvAOHh2oE0DFTlpM4izyP0+gGpCSWaiLCWg
WGEgmEdehQmXVj2Xaksbc1F7e5/pnZI+5L5vI5w8aSJdC9TtEWVUHa3ni5EDOUX67S2uAagwKvw4
9PjgTD9Szbw3Afh1nlO1h+dFcauW3DO6zOuR7F6Keh4kIf/ngs8fUKObpjrTWlb9URy7BH/Qtj2z
I/NhWtXPp02qMiDntoK2D7tNL9dHXjmyLYZFU00/zNzxWCFoW/lVis103afXiBilWZO6vQvGbDGG
KqofZVCXmqTHJ+UHOHRpZ8gMTgcHv6hMAOgeofSTbo2Z6Tpbh4i15qya0HIfjmWtW+aDmvPTy1xb
vqBl0RDHvYiMOfCthH3qSBIiRYQynbJe5KCVj8y6dWq8ImuGQdOCYuYsJXeRrSABztXvlQScgM5F
PUI/RV6hmsjvuCUXOgpyEKAngaGSQayaDnzZ29phjKagxfxyBfLrhGK71V/3AxW/JrGyi6ihEqcP
8JdbLkQw1VCwrzltI45YIjnXxqvG0NRMXnvKt95Lqly+Dng8vh9pdtz8gtWCzKJq4XeT3lmz3A0f
kFYOtOK7MtT2ZtlddJ1oGkFvMubRxFL+vrSScgZYYDU8bOetWaDqmLhjyz9d9gZDkXyuuu6+/6/8
KE5SV2jt+DkmwBBgYlO52P4Yy81AyzWOcmYIVQZYiy4XfUr9BZ67/re0+fYieVJoA1gBbL7EWwnJ
BzocE5bnuBR7oSG7Ar3AqS3d4zCJlDK0NVyaHMuz/V6Y+KqTOhZaazU9+P1cRgYiMbS9lIwoj3Ip
ga36tXs6ZCp29L4tsENgKQzp3tI/xUyuruVhwY/FujOft/AQjl6Ai+twri6lHzxdfpC0/qj1Hkwy
Z666bbcGhIkA8G4do8r4cvlx3elGhg5pB5WBo3E/87fao10J3mdUBaXvB75BCYkMJSMjgXP5e3lM
xdcBU6DXPZ6eIzg6F5zEaL1a6PBbR39t5c4TR0rueONkxRmt/Ya8RF3G93JpHiQg1ryW8CiTvYMA
tT8+GSFm8rZL5w+Sx6vUTYUaCoxWNj+VEb+fZU7yyjcpum9CF34pfHJ1ywZtDwvSYxQDR13zGZi+
JDHrspEifc2OvvfN5TMyTIVECcpoq91p83bhVOQcVePCAvGPxMMb2/32Df4MayXOzvL6kYLv/Snc
WBaoC6MVyne7LIILj0rX1p3sPLGsJfliFCfypUS6TwFoBbc+UwABF0uoXqr3BJCP3BVMt++bHHLN
mZIm75Y+89fQBUPYosEfAt93naMbaYf3xQ696GR7HBaQFqoxQX2upBKi9n6ja1Z4fkVIjll4/jVy
+zezd+9eRUU7IOnBLgyTON25ShI7RHq6WwcSiFgNzkFqkdT2cFD+IWdfe0VFhc3har24OKT4F2/n
vrhTKTG6LsIBD4p34c1uWX+5U475oP93PHKMJ78zt0biAiHK7m27KCr8qOnRNyaLsMuGQYiWya4k
c63iRFT7STuYA7YfVM2BVZw7l16OlFjNrqW/iq5GqH5AwKNYjv0O8KAk0wLViyJ0IDQ/QCiGpz41
bGipoexppCPEdZ98mJ8R2CrbQVeP+kTFcRDyAwwkVxnm7HGhC2AV2FCZIgMtnGvvlhj+BsqIFev5
ifCgRFY83mvCl7SkfF+O3r4lcDOhf5JjU565PzteHDKGUw+Z7uxg3u6DBGBAo6CUJmkDnfye3t/3
tRmnNKo3d1xu3xFtE2gPebvTjXVKwXYv+qvP7FhNfrt8sBFBc6MKZwDbZYOWAaAR3GvYbVFpDW6W
oiYaAsodGLHWaWPbo46Str672uKJ3aPGE0MZJYTRx5ZJcqOlkWCZZab0cQ+4olIhDe4kj7twtIo0
qL5YWVaPhnQHuLw0h/EH9lEHwJ2SD5pJJKf7M5MSSSWvtEk9DJyf/H4JVezgm44sZ/wnmNbp3qTp
h+g9DJPI73qMqXdf+h0jz4FY+VgmuAZERFXfsjL50e3TNp2JKt/OxFM0X50PXI/bk03FPbhCy0+j
GZ2hfHtL3N6yGtt8T4am/OXfcRwWMU00jl8Ev5K34au3tR9V/muzbEQuhSThF0elx1mp5Jm9phbh
CJhGf3wfK98wbHhvecI3A0o3jZfnljwJYHL1BsEsZvPktrny+cKOmwhhTKc7sxUxeaqo5qOJEF29
zi5UsElkcESO7/W56HYlIXWBFWu0OY9TlG+cw5jSdnBg8RrWR2FqhbimUbU3tsYMqr03lsRI6OMF
TXda2Xd9oMC4QPtZLwWXGSwlk6TH+O4Cf1PHQrcINzN7HvCzjpyIAh2aQwFOiGdI7W7YQ3nwrC3W
EiWDd4K2eAQwTgpG856HKcr3FKjJU3qKo09lsgzNOgXN+u/7LXWyggwwCPyHHbh+t6EX7jdIoUYU
4y/xcBxkPYoUQLN8m3D8/vyLkU9PoWNlCgEkx+BXw8qJP86rYpd0d+GnVnm02aCy58FgLLdA73Lk
FJVPFm2jlXzdqjq1/1YdqDM8iRS0Ut0WcOMIfAPOEZnPQy3GXoadyth10GV/DZLmhM9QXZWx89Z0
JjV71fmC1xqyohrLSf9UeDiOSG7NOVatV9/BW0q2SmFpVR3WdGsKrkSieA+foxZ6FpFOnFqk+MW9
6hZ9ybe2kpJhiyAWgnabqjHb6I5y8N02CwEMnUSGnga+Tkr24ncNDUVT1t/E+R5P+teJ1B0YxMHI
Tw8aP0BipSh88NF89a0cho/xpFJlpW1QfBwCv60IQW18LHkS/cN0P+W56PZYkD/HJv5FD4nt3j7u
Se4qD6JhlDy/W2/wrUIqxmMddEcJuAmokkeA1wJ+P3y6iIPRSfp1+fawH0zCKzM38Q6kO+2EPHDq
nNNyo8+7TKKG61gppJYUiTrgdOwCEyG4ilC9KQy6ICIZitZp2lOJlTCupscwNBr9sGizKcnTN70f
48tZl0VEZ3edDLzdn3G+0PsY2VqxreZNMswYSI26F30zafJydYJJ+IZi9/iZICl9Z6V+oitrWBRp
RE9u6K76/6nswagHiyqt7wWKwlkRqPSjzLME8q1iGikayBAY55teaNmBN8+cNaDWDvVKQ9t6dVtw
Nvcww335GjX6f50/whOwyyqHjCi6KM+zl0jzFvIwPCfOhiliD5QwzvXkQ2Q2C++u5ayH1Fj6rr5X
ViUuuZM4NAOPfbIIuN2ecZXN5Pu0DZNCc33c1mPDePSm3b5rZdtUEWA9sOyG0ZZSx065/QEvGMiK
48E7BzP8Btkkp1zEnPF4PvabzO/SI8hEnPAropgpMUqbEde3uFGeRgljup54dgeN5T7ZEWB9m4mr
YGpzKku4IRetj2EVfSLo1QiYkTb52T2RUu65q4uBOsl+IsyDfIstM+O/gCaeZkJN04JyqIZOvt+r
L1Nm5/gEQOFwNoVTthHxSo0woQuqxcFyNL+YtiUIvRx+gaLEbeonggUPUUacsbHlBrRFtuMPSnMu
u74oJzjA7PE8L5v1FWfo7skQrFjRjQmGOfqhzghKZ/psYzIhqwev87FZFe74QhJs7fedFjAOVedG
+F7YNMaDn5TGjtrO0OOZeTXwrCDt9XRulOxf8T5a2CtdcyDiaG+GBfpBYojhkFjMgkIVk2p69bz2
7exJSmik/8zXRcjWL3e79Num0CsZNpt/RMYFDezQNRjKDmCjzQIO5hiId68Jg8JE9EBXBxeXKK6w
xHZdDRLLc/+giQ6dCbBPyHyLmnhPsK1Zj9wc5P963AJLOd19W4wwdIJcOhblGnxf4s2az2a/rDU0
Xey4sqbAu8a34XqMnE/fRlv1a6NKcMeO6t9KKsTYi3E8S8hSh16EX+E/dc+5yA6Oyz5lmzg6VSXQ
VrK8LsOkpZ45sueM+cDDLX717RAfGfF313o/H+zF0yv8KZNxVmbJC/IuCo8ESPgeuxJzYSYUZgDR
E+FrCgVzXYe7tHTWTnB6qD+bfXKN9Cbi8IBnH8ZcUnILXXLElcvTnurGh3SoKTZ1J7u+mUzk7dPp
1qh9e/6gLk7UKItLHBBIlfLwJmBdafv6KXdXre/g3oA/d2PPcjzEy869XGVIVq1axJ5W0K5+mgpL
+aaB67rLBp9+RCTK//x0rejOTeve477KqfzNqzY8W6EdTQG/L/zktVYusHBV+AN7AaNkXCf5qsPX
we5b/DSCiE34+BshrUobkDOsiva8/Yb8UZP3+vKps3PfZbAeDC+plu9sofHdLr4hzM53QlCvwNMy
oaAx0VWxnXmPNqgkj2DIsQBiiyhs3FCvUOw8eRrz/F+H2lPubIr1I/XgwibmIivKF+tAu7okAZAx
zdfrTMhLcTXFpV7zWubkE0U9vya/scusHG+SrKy//Z2+d3lI1niPMvfg5RQpNE/2mrr2T5J3XjpK
mWYa22LOZp/uLrDXrbzMEcBSDsGLWhoPW/KZDrrjgAPpB5z16oQ0N7sISUk3Vb6LBgOeDStsmNkr
f88XUNRYPhyTjC2+BRqErMNxWaAlCp6zUnnysebiVKdKE8TOkERtjG3kjR5ncNAvoZfO2Vpa8Zoa
8f1Mx8dmz0K/dg4D2RSt4ZOG5utEO9YcJxwuQAzC3YWmo3FPatZF/5h26W4dTfzcyRCbpcswBrh+
ZclitWv33PmyoXWwzo8wo42zTWDHCrUHV2yDnvnRlMStv8ISUCfhBad2pYsep65RFLhoCdN/Znot
NuXAQIzvyPfTdrw3EL9TXJLlQZFt0n9DlJFP8LAgwul8ixmT7yWPJ+HrAeQrttSOfXxoLAf102DP
v8z11RTqi22WtgU8qReZjiZrix09EN47q8U0Tl10U+aYLFU0cYIZEc0L3C67XPxKFiqvoeY7yOAn
p17v4UBvkNO4cQ7Wo6gbrhdPKdNkaCSKwcCtVZ1Hbbbty9hUY9/QdBnvO8XaLOrIjuz9AHQ9W9S9
2URZAKx/b3/+ouSzf8AECz8Z7/+WbTYOz+hlhzi3A8fdWbqfFcSfuE8AlNLk9V6zlzaXr3YQ2Gn9
kAeq6dDQW1jUTO0suldA2FAc7sehO1DCb95RSmyVXEUcH5st+Yxm12hIP/VlDZOA0L/j666wjHJN
Gq3d+ip70UyAD8Ya8IKu4veGrl/YIIexlzKanzqSWh9duZocqa8Yh6ZVLjpR166hu83WD3NBuGlz
Ztzqd9nNtEZS5vWGNRzgJuyPoz/aNR/dEJOoQVmA57YBt4fnfgsoqWXzT2cmIiIaGuXFT3d+0FUo
dEswCq1oSulJn6TDhaJdBfBVX/j6ndMWX4gFVWLekCSPBcSuHLPho0myO2QDz24yaE9xQ0Z90pG5
S1C56QWtNmLXWuj2b0nCT7q9O8HOiyJbBJCxvQlFwzk/680ofXnDkuC0psr+BhbDOyVye+hQw6Uv
oxIMAiQul5y5rkopfUD0t15GlGyLqJleONkCmF+fPLXNfewFaN5/w268H/lao33r0GexIJUR2WhB
1dLJ7VaA3Nx1rC1GAOH0lwCHFLBwdLFsigqP2MkheJhA/TICLDExBowfFt4KvhTTRd46y9qX5Tk5
rySo3xXPTCJlfXJGTNHT8U8aN7wz5c3U0Irea/UVvHIA3vGsBjsvYrbKSFe0rLQ7qE/pgmgZbNdp
anlAOLShLTSxBvTJgDaXqiUMeYvGbaxEnIiXjBoC2o1h+QI+a4LEscQJHRffB4NFOYvfQc7MioFw
pLrQ+/ReSIbfEtMfz26Zb2/kItjgeXzTTAxS0d1lHEvrYCNroYz99evIktN6LHo5ztHiZnG/A/gM
/FIbqJAcKLVSZmnUFyuX+7jMsT6wAExt1tgzPXhT30OEzBsEJABl1m0VJ0vxpw87dglI7bCxvu4h
Ex56TnxFGLzksCmJnuABr3hBqpiAcIszOG8UaBm9P8Hh+pNq3rnBvYzVctSqgfmbsEWEVPYgb14S
DuVKgdRmr3KIjz8okTj5+uKGGIv2cdiN5K8w25KFJqxR8Kd9cVSBG21LGjzsAg2Q8oKYvs0JRF+B
f45vd6pTFkTU5NVQ8PPKkxxDr9/IjoNYsg1liuzHQCM3kAgPcvjFHnVEd84+JqOv3rYnaFNEFrV7
aHHWtzR/1OShdQYm/nDgoXFtL25kJh8AzZv2xyL72JFXVYfUGunh0OL3LyMoYMBfAaj05HC7E/Cd
UZEqKVMk27hxDd75wXib3hHCcBPkIEdAHLwgWwnEIOmWB1hryxxliZJDsUQb7xvO66zTyKK6MqqJ
UIURbosZigL63D115qMnPxkTuGolrAgHXUn1E6pv5OYyIOEW3C5YUcDa/9zCKfrMhviObVATMkyt
COyXNf6GUFzryLZygSdzUYkS9Ae2JhOs6THav1p60oelfXBLLKCfLck60mkk/jBx1KswZ16OjoxA
gPRNXRA01PWT3mzxD5ZtpLJJmgbBjmFj0hx+BG7KO6XPQ0UeGau3f3xOIh48lBeujDx04FI50Aka
l/8nOHQaYItAKpW5QR5cjkGkkKw35tJygIcKQLGiyrBPxkZL6EE/cJeu+oS/IHuul75cXUH/hStj
1ot5FxRkXGAgpLMjeLy8xCLOoMBjVkP5T1zbn9lGWu2pJNyQWNX96F5tJ+wbd1ETUaGax9imyac2
6Vi3vR6C+VGwEysMUctOKyo8nwG9PnpNiduEXMTL6NsFRXLGSLERwyvlA+dkhPWhLKhVSfcsqTa3
wOWDku5xuojEyEaimLKO3ieQJGREZrPijGEg1m20WIgkCu/o7+4N2y4ZLgXmBolhwm7JbEv8uss6
TVoBIV+HZ7heRpBnT2ToXvSXsOk/v2EeM+mnIzj9f6bmB5ZSIra0dOZuUTbM5IsJzMYBcx0eYfpL
I8cqmXHO5zyHmAd4aAkMCoAdnp+IBa/DrEn60yp7rbdgSku8/Yg386k6ckR9e5B8N3VObELkLlQS
278mfTjDVM1kPSg4kHXcuka/74KUEt5ly+A2TwXKQ+hVu8D+t0ECdVWXOAAOR/JMbawJTWSWKsK6
N8xgDVX7ht299efgS8SZeGBTK+W0BW5Jr86hm+DAWZfpB1GdobrGuRcfUNEeVN+5D8pi4O/vlT0d
AgJO7DWWCY1PqpVdMRSjikkpcUzw196059mr+j33s+bv0fuVMi006ImgcNgrvxOtIBAw+9EOOudI
WE9GBRfMOXtSETBGm1kmPT00n7rC8iHAb5LkdoEhjX3Vx9ay8c5tLG/0jP4h4Q27P/sgFpS7SyAM
7MIr/cfp6hGhsNWkX8qhuEpZ3qjtSzrnwv5pNcCx6T85LTHf1rRyGM8MuHBRV3NenxZ4m7RbgWx1
RcB4nPbV+KGkfJo/krhdozEuAcvQ1HpmJCDiFhRDjTYyvzQWjAl4khad3XGPM7nPownjeT74Wwm7
UYpLNFCo8xnCMKy9IONboYKSevTWKLAWoSZdFTabcAKXVo7ZZph1MORaphvA2XybNYaB2KK5ui7i
mgldoaJtRQMSOJ045cMNkGFfvcXlOU7wSTnGWgRBBI8CB9GT9RfEzVbhJc0TfBIEwYIcJqb+cvNN
DTxB/Uy6lkMDLZKypUdhKy+imeH8JsogndaQCCT5eVsB6aUp8lo87fmZVdE8iEFVzemyObt9SDyA
fWScllNe+5COUg+rFXimg7cOS6gPchhgIGKtlG34TRDb3OIVuYjqAOGmfeNe/4sOTBZX4tvld7D9
sbTZi0H7RPsQo0R9KhIydBmk78lP2w4v6b10AAAiK4zcKFbzDrLOo77K4q5lEmuWYZAH9PQMMmWK
S7Iy/aV2sVtWZ77tHDG4xJ7LpsPjtBSstnlzKvSl0xj1Tm30xuNtnqhfkprmcF5iSKkjcYw+//3/
cHSXrw/3Lx0yxbfhJoQc+1+YsBVs3AvjGcdvsPC1wIBeN+BGqo7PHbqM8V90Ib9mX4ytpKPZAPel
u1HVrhr+AE8qWpTvbOV8bG/zTR1OZbld2YHieAFZ5GfML/yCSiqmQRTbmfRltogMMxjpnsTPe8YA
MaShb/ZnH0blZiwAy2iVL7ZW2U8WtJ6MwSWKE+8UFy3wmPTi31jA+t0XUJKrcQoqwgFntybX8woc
uU6DFHtA+hrbeaRTnXyrm33DjkEy+A367DTJOeil97ArZwB+dEtVqQhVt7QpDcn1hxF8Eoe8VG6o
dB891NmhlsFBH16z4jNTwP1IAZg/VHJqmRM/Niq/qmxqf3HSz6Fq70FmvuvipX+I9vvd7ZluwNhW
1IL6QcZNUyWtyhNYdVKff8Os4pbyf3/dTFiBoIMO2MscGCRLCJjmibckxBAUgFFB+zUxgH1iPiq2
+ztRkLfQi3zzydTpLQd8aEthUbyArBeFx9lvS0Qa22680dfwisjpDMnTF+IbM0l6CCXMiAvOlx6V
jYwDA86PcYiuF8YdbDXI485u21KNRFrj7glkdLbjm4H2jxSukQsCtDJ3OLw3IS9ag4plk77CZyt/
WDuCDU/eNxPl5B6TaTxiGWgBaMGKCiUVfLl6fAGaPTS7yJgo7kSMyN+hBBSaIBo44Awwrmt/eaiP
XWzfEbdU815HN9meeDbo7HxT6Ro/Xu2BTyV8/hQODkFGRyVy9ANh9JsMjJmbjiHb+fF6R/J2VS/D
DFT/p58NIx9V3P5HrWbo5szrUEw4mpC5HR1zhjK+LcX3ise2ZUQZlNEXMOsHcBpyvGnJxqVaI78t
6PyMbvNruU4WDU+4wVdJwRwHlFJxsGiuiFRXxcNNryy1+YpNn6jBhGS2G+AWaH1s6uGLMSMktYvw
YZGTx6Vcs4TpXrkbR6Z8mDnhW9PmfuLGzV/BpZaJLwRE1mpmmvS8gHpl7obd6LBBPw3YlMXnkwhO
+iM1FCgqx5wtCDtp82qQq2ax23lhbJDC5WH78WGqNJDz9A7LWdPQXk5eGrW5v6rJp2zJPPF3WBOs
KxO8bFmvJdKRD+TNDBSckDvjk7OHig6LoYUCKJLVu7iCFdTriz9tm3hW7vY/72DzgxcbBOtoIhMX
hilOXEu5Xqqz8Uv2FF7W51fBj5KzugXMg0oPL0xxVw3qrKKn0kWZOh/OGQc0y4HTw7BpoJyFbzab
gsDBqdqJWE6sIuGnS0wlKoqYECy5VdiL6gXEWDBoK9nJOt9kiW86yx+RPrFNxrn5U1XGQtCE5Tpa
6DrLzu+kayXaBZdf3t13tQfWN71dsm0LM1ehDJ1S8Dx9fYrVSTW0j2kJBZobXD3+TdclSaR4UQ3/
BfxJTPDkRTJe9vQ9PkfgBgM/JGGhUDsH194xf5YNVfDX8LsOJKqUGE1ZdvOMrOBB+gp0pXWtLvVX
iPUaMAxnLTI3o1M+ULDfXDxOqOC997AT57yAcdqYXzjDge30zMhDZh0VLWpMvja/th33qNl4AlP6
Mp+ioY7/J1ad7gBmg3Tx5Xqe7zwEuCRi10pFdVjvjkJnH0fU2fmfXE5c1j/ZBzbbQqMj20pKK4dx
ISNFGyAcisCB8fmS+4CZ7b+4OYkxB8iktzUnX8cQFT9t1iI7JuGSceFyfUo+zHWIpvHEgkArw26i
g7fR3/T+gZc/DN9n0IcETr+CNyohzxxKhhHHd1GNs6N38mqnvxqhv9ueb/50/w3P+v1hc7RAwlwn
0xQqNXtNETQiGRoY1FSFTid6zO/p62Nqb4Rvb8XA9TiAJx3aA/omx8VG/ofPCnP45IDkVJykz5io
iKGtCLdPC5gNJutRbXTsURdq8X19gMy71y72w7nnZHoqKBxUaygpkB+ySi+1KEsHINVWnNyiDvEd
awsxfm5bvnBWN0wmsAIugYN6eB4+IVgrnT1/WmsVoOma9IWLLhhLPk1jEb0QZsV5Qravvx9/O6VK
h8YvXlCZVmw4Beldw8TGalWQWBML7Ym9dj4VmPhSm2LV70oM8XpaJLrBvSmldMKlgxwGl+JS4Yf8
GwJ7CaXuII7cfr9/oSB/lsEyROiSEPAbpMS/C9K+VsiMJYcq9t1ADpumYhCxtk0Ox8BIjtba704T
Jx4pd8gyDxdxrYR5vKEbGvKoOVlqBfOT8XXaGlvPy6XHStC/EAzF+5M6quqlYczHtdANLBtVFi7w
fQXUCnkbXPNEQ7NNBwFhA8TBh4ZtZc0J2Fy3tITIKSLrN+v0vn1JSdN5Wl0KxymWBsvt//W26PlR
6Cyh0AtRighp49EnmEqP0foxAXlSes23S4VQzkaGMcdEAqY5qo5efJjjdAWu1It08mlXof1mWt0G
6FKtZze/yJ8RFspOBz4KEZhfBPAKsKhxO+tFsstOlQK0rE/cA71l+p5IQL0AvG6z7ujtpaz4lYIz
SnOF+Uf7lnN5axdecBIailOhVDW24K3D64QOHTdfb+0v94Gg8v+D6wkdu18ar5Gn4j5/TzUvKf2+
PdJhaSPLELFtVquy89h3lkY5AcIQqJv+ZCm0MIJ3GTqMUvQqoB0dOydHgHcKKLL4GPFSG6edsTor
1dn6ZxiFN+VXhrOp0X+0TTZQHzPJVP1vkpuA9zWXiqgGDsm71p/kpxqX/yyCLAAnpb+wIUhmDP8H
Er8sIK/i+lOAEaU5CQn9BIMLR7FvHgT358M7aKIvlnSxaL9nStT+DxsDW3jAKvOyAqF04Xbr2idU
RUUrUjSw0Jnb/saIDkp1vBqQ6MQotFDqaV4iZxU8oivOeHw7cuIC+TfnRhLwTAFH3zEy5XuDaxBx
yJ+p5Bldn4LPzy0oSxpPzr9MeGzTIzOFiifCmDbjlxOY7iqezHjJ4n0IrdePtEkDGMiNszBjpqxP
cP7MqvkFc+KkG4sOEnmJW/g4AI6lmPorwUBcO34kzVnAS2O16euIS64z2g7rCg7fBYyYoyzzfOD/
z53zIfBrUniMhJ2BIt88lJpYBN9QoSihlXQXVctLbbPiRejIVPbv7FxPIO+knHt1Ex+upqiTBn6H
YPTKEyqZmGQwDv1z821JQGstu0+n/wFPR+FR1axRJ3WVhtMTTiItOh/9f/XKvUaFKQFcLI6hEpTA
66upmDi8FunlPNSOCFVQvtY4NKrwY19qXKIRpB0PyX15mzS06FGthKM4nTyiysPMNv+o8sZatG4m
RKYceewarCaNf5DJp/uUwngtSDApToLBW0wxzeHup6hFDw2PwSbnYdIctPq/HCFPk4422EHgsdb1
vZs/KqnHw1HJ+328vCbSxOt54ljGTBuKohMMVn1IuJC7fWC/GcuZTTGUV5l+G5mmGw1E0ZQd3g3e
zl+f6ok4o3VHruIuTUzVGdlnes2AoAUOwc/FfHAHVi6tEWV6p0BrfJdsmohZIdd0oc2pZIsV9XIO
LOnHkYa3rz+nydx/t7c9UPpV3EJmSe25lLp0deC9fUQFUwLtQHZH7xrFGI9WbzhZmsBEj756uEfo
zG7QylAVBotWsmXt1sXVRYQ2g2vjqqFEIlrjyd8b4sXRr1E/r0NtQhWlDHp6ubrYmQ5qVTk6dRo9
cA0IQkP4yQyYsRRqKJdi5jMkDp2S+5iRoAXB3ZrE2YAV9kQK49/+bo2OcFNUZvF0Ht3zY9GkX/GJ
COOc2P22ZS0zLVYzUDyiPGETx9wsMgVjGcoJlWb3smXmW9lhUy1Oqb036kS7Qz5bwjdIsm5/qUh7
6DKBqyGgeKtfzM28K0e9Xas5sWHzqt2dhPFKl9ZdvLlEpu13Vx5SS48RPVJ9wFVHo05iQRGWksG+
Bsg2tl5nAEG+wxaFFM/PBD+EoUdhGgxYqD4zOEJLAY5u6K+XoJ+vUCE1n0i11rwnTEnj+H3k4eiu
HQtpu/Z2rSqSVD15NWuY5nPK4BO7APA5wjRdvekWvf4jBnDcUDMyujUNHYqVZ+kviQgoTl+o4cWW
5m6uvpnxI8CNnDCkdYWeBLrqVnUw6YFsohkK68bi0nOpD/SKmhXj0sg7n7C9JInjwVgNkgmITtol
qPJUp3WZjQsrZ5rPrdyYPrFYbg8zhpyEH3bAY0q74KFSrDOxjdBdKXCqR148FmEcwJ0/Xs6y22cj
nP5th4PQWsqluIZ13dLxwkvWocA9+h7DE5L1Tq0+g4bai0FLW47yRC9NOBO7GRaY1NpCoWSawcy+
Q77lDxrx3q/LBhY1Cq78CvTQ6gR7XwIBUVfEikcI8u7E8dnoA0LqgZQMpEhnfDhMS8hVFyNpctW7
Yo2dZ0OBGD/YwvR/99SA9E5aW199xxK/y3mgKCFyqVLzdP0ylwy9I0v9uEBKXbQzMPiZRaY1kW25
6w5jF5ZN3Ay4+GJbpfw/Px+IRSxEgGsXWeDUMsSvCIqT8ASmymgVkWusUvfKrEdqvbqOPOf770Fl
FthM3sHBNcWlZM1IZAR+jujbpe8Vxt9PQVMJJE+hNe6ovZYR2nS8eWCrQL0/dKIoGqmNNjI77yzD
dVoAKK52QWWdOsLV3NqwkjWya3vjVADdZ4QBa0RjDOUPiwN59yK3cE2JQZi0ByjKBTBNPKlzbdYI
6s6uMQixD7jN9nzy4f1z7ZsWd0Zk+RDGg+xQkf3CxESKdhrc7QxAqgtNQNqvsmsSkDmw/qpo687T
91oh0tZZvZIt5KQ2edTv9DoLXeJw/NNQSy2xDWEEHB/m+HalGjNH+Md4GL11ZHcB4Y2GDn43X4k9
ZNvQS2CrdqSBlYe1+UWaW0vbgaM5uOYgUBK1uJDasuXHqVZUGZPdjKy/VYX1DNSM90SGf0U8OEXe
7GiV5edOlvMExLk5/go258RtvS5TZr0VuSdqBNNhnLAtJyWPPokvmnIfCfsQIUgCY+nfzCWrJBSv
3mE/b5NgNyxW/mOrbswMB/tdBq84tCBjyocjoT7GuZnpWSKzajdFqVLTd6MBQES7V93HSkZA8kWe
oL2AOec8u7Q6NrWo0ZWL3s1Bje6vrm0KKzsjglA5CJRwf9NLMlM0F5FFC74+8hxjXRORMVozcEgj
zSOPVjFJvAS+MiXjKNSuF8i8waaQDdvgixceGAspvnxpW/TpFJ44US6NhDZZe00xXoNnyD/9xHkO
DRnTmTMHsdzqhfZbQmGwyBZPZo1z7oYA1g4+dxdtCqTu3I0A2RB9rbhuSoqDcjnJKsDkyCB1tvgI
vR8AJ7yJ5AZLVTmLqvHbkDn+CYGHbPO8E9GHV6Ue02TPG4V1Ht/wPjjpzYC4DOrNTSOWx/cDpa2s
rsBNfTqSZbxZV1yThurnX7WWJHlAiCHNWz+4x1AgSB6lRXknsrYegQ946xzobRIdvwoNq/ZQ8XMf
36gI7QvqRobYev9eB2JvcWp5EM/n0/N+75s7PF6I7o0RxHDVPmkolEsOAQKapkH82eL6DoNCr2dD
DoxjCQEwAzaH9nqLv8tcuuonRfA0VC3KItJ42x/eypAQ5cJawa6ItzVkKiJ4PE+MDZoqwMbeajsQ
Ue4ZRxLUPQJzxUmwIitU/jq/wz2nEqZwCcpknN8fGyRaDuC/0dt64bC6azJiz5OSCvQ75qAWNzNw
RtJe3Vpm9gMytcFYMun9fq5edjCuPgPHQGpw3jT35GVel/+fhGLNgkjQ3foi11AN0kHqLkszBb2+
P/u3pwH0l9HvLXYv+E2idlx/7smo1G06eeKYCFdRv/UyMo7DZwZu0jD2kYh4ksDNIyQj3a9g1/47
FvKeUpWNoTDcPYIW4amFxHkt4nZyokW8M1bYRnRLcv3gls1e+ie0IYQagBomGq/Rr7Xwitkj+Vmb
e3T8Bgdj7Oo+Joih+CngLCfAaRHfqINO3gcLmsugL8KCv1M3atjSWQcxDp0UaV81RBdwbwZsYmPB
YyboOsNWaOfJyAYwb17TVqXIH3DD4HwIKAotc2bHKUSEBlTTFEKWaZU0JW4xqqdchJ5/3ZUNxgjY
NH2OZz3Qau54UztF4f4oND7CaVrbXNx+107aHEO+rQmPGC2puDrI5iTVcEjMI3mpz/obdzlEKJwd
fEVqEJArWFLp2u+IRchaAqp1mIIeVfdVxWLtyXOwwZr1C2RmRtyn/95OGVDc824vqdm9jWhL4Xxe
2pFC6OoX4OHrv+YQHDT5vgmpRsrEjO24WfpIQ/HYCvPvPlZxFskM+h1MPaZIzdWK2qqOixKGKume
Fi5ltuGMhmrFkhI4heSk6hLDfqEQQi8crBq1onTfkqJZS5UyXPcWcVmzTqg6RrVoeSjTMKphaG9x
nwzllI7cZ6kCXFxUzvCF+901oSX1D2e1V7YV9LsqANCH/wx0Ef4FA47NhMzIbdOd/6/ReJJiiNWM
oCMCHgmhBOytJfavNqMwu4PofmoApXKJ8oqMRFqu7fYy6p5c+Xx0xMW+X6Ve7UH5pX8D3zM2dX2V
pGRWs/f0PagLlGpTOmbHBi/a9TGe/6B0wzrMrybDgScYCe5nAVCDcDVAz+pYs0A6yAtAegUEc2dm
pOkdWTFTCBIwTQAAWjNRX2xad1p0jo5AXhbA3GXXajQFehdSwyZGN+nkensXv1S/itVGC3FDgEhk
bciGGAFD/hNgEoH0QDTft23N53AlR+HmnYCznxiRgk5jHJViaFW4Rrs8phmIyPu1sAVffjzzBxro
xkiImQTQ3ceShE489uV28vitKBhKk5LbSPgNZrjAXGJ9Dz+lIcXP11xbb3VHHJeCDb4hHLTwE1lL
1X2MmRO3LDy9VAIlW/Irg0ZtUob2sgyCAn3x6g2n1pfYXa84lCYDP6sDBYHKtHlkYAmqcLIvLBCc
62vQBB49/UvIoRzQ7hR3yqBBwYClQoj6tuqU40PZkA4dsehVNd3xbXx6da/sQJqBgLX0jjxJ70vp
Z6O8hb/AswKvshd7wZ6lvWwv3v2UMPcxVD03oo5wgOcPaFGo6bNMJExTvKeSBIUA4LZfoDS40/5B
RsJlAtovlRXLhGD4cSOjIwPpcThGECw7jTGX2zj0fqvRwWRWjbvCQnlPCwcXEtAFzwX4pD54GYuY
uqkpYhKnrKQnfBvRfZlsPgec6+douDtta+HPPM70zmgOmDyaMtYHpqaVnkr03qG7MFFbmmHisN0N
+jqwbV3Wi1+bABiXYKddEktbqVdJuQPdMpvbOYW7iGAOXort+ENzJllTrytZ64HGW5KEvNcf+6zQ
/B9RRFPgqS/4tTLgXgbeOL4+hd3y43Gr3x4yUReMZvPkmn5tr6UPJIZAyaA2AT7v0kANCzUgcu/m
E22/c6dfT0PdG2KGdMmBEv7gWEAMUQmq+c1YTDWo3XiaWi9bn8cV6+Gqk6uA56VpuW6Q+VOenpq3
SWAtDSGcLVEoPOBnlWyp93sPKXUZNpHGXX53qqInoqa3cEsVw5d/ob/hFL3Z2Jo9q/eJVJRhJY5v
lgZvNSe95on030aMNMDU0UhZcmAcGhV0NOnrDSJet2GPzAyDa5NlCYsU2+bH0AT1VUussrGeVMjm
FKRjk/h6NMGW2yAcCm7Ayv6wR8Diey4wsFfnJtB8ZsjcVIWYX9kk98JAR8QtDVKwU6eKClAfO9rX
1AxOXckGhWIoQA6y5TI0HRhO00HVO1QCJ4Pgh0busme9Aoy4V867x33f2Im59ekYtgmblafZ3pCO
IDsxKs+NGzn4JNMqtlpDUHgx3u7dPLk7HtPMdRAHjPTb8kof8sxCJpxgAy8FcgK/uIq+1Z4OrXhw
aRae9QCGoPwp3Qq2lEGeB6CZZp50xcl5e615I+DUKYGRDCDKnXKHAOGixHphqM5LTi52jPTOeY5k
O2NZ1heC8izxwnhiFLNviVqbn7kbCIcvA6b51m35P5LMyRiwXyy6N8vJAK/Z7q6RlI1/OMVnTOxv
keqqbiMcEOZsWVUrCmvN8zIrLqm6WpIh0A0ZokmiDWRk4wKTbTlQ8acpC+8D17ZN2xEWQPIRWend
YtqRVqHxojLYe/PmMLfmU245rhi+xiiYmHSMtf/gV+/HH/j3oQTeOx0C0AJdDXAi4DNvxkFHzWke
EZSlGyV9ZbvP1AuCb1vBsIQ1bvFaeSs8ud822LHwhvej7aOQjEgsh31B3jVd+25vzvQ1ULKPrBL3
ZHS28S1LMu9RGZZbDmyAxJC/gfY4otv9qYaEvKiiiHS5taizcrI8hF+Oob6Dk8Tds3pUgsAyxSpO
0UpWMTnpcYJ/FiFP/8UPNd3jOGcFlusGdH0/yJXTjak8DnaAn7IebHe+hyVwNdCgyJuSbsakUNqF
mjWhj5px3JDrEYSnT5yWNOcsmzgEiqaO7ucxLeT+a41UIANa45TZ0M89Opv7TWKH0eOJWRcWMvsN
4d1vDNvOHWeC0sE5uSWpLcsmiMKh1y/EyN00jtqCxpmGHyMKoCInH0q4JYyJUIG+2JVCHNxDyuOq
LAcpJ8AVbmfQxZDkr+1pBhDhvf1FV2SNzG4X9ieRgBh+ee4NFvKiv9Z09j2A1+9ZrDjc7slSaupo
JIaaGh3K7KNuu5hFvOmaiBipHkadHrTUUOvWnyBOrB5EwckJmwDreFGdv2r+vOD9I3MsqpIRNycU
+xt73vIiWMRYUFNDiYtG2BT0BvgpLrcJoaVg4XQswsyt3jXlxu25C5vM1sZ3BcN42jbKH0QepAVO
qLAfXk/saWhBCSEYEzhw/AAwmQmN4KBYTNwWTg48K4Loh0bmEfkO1YfoaehnWHnzr2pT5QUTLAyq
AgT0hL7mg6kQEfCCNsNSt3+uC8tOaSvr61el/fsvji4mOf0yTjgHabx9X47Y1ZLEhZyZydaSl5L9
hiOUEu3Q8AKniJAFiNOqOiFLYJsBgnW7X3/v+iqt2TywETFl/W97As0AxjOcnM0fxibDXJ78390O
n5RO2Gy42kWBz1cyDzFzU9wzzNdFTlQtNzXgDy8YW9S4E94jhv1dHJBVv/ChomQloSgIisA114U9
5TQocpAA/WdrU6MmTuOa6Emn2oGr43MVdlstnuUdbj8O6WEzmzPfaPl/dXmJN/0ul9uOfEdYFiC/
t/uvkT5r66U5dx0pdW5hRGl+hR8IjpYlO5xaoREX2Imr9fLeZ5Hiadlsu7St9g5v4Dy5SSiwhBUa
YJZAh8gHE25MGLVlcyOTHmNkWlbHm2ta0CFSbMEUbb495OYFJc5Rqamtx1k4N1VWr748emAYczZl
PfVs9RhYF7a6uKEb1XD4pGAsRT6HdKVtSREAqJ1tXPXzyV0PQ42hvpPHmJur5/o5EV7c15/hrL0H
bEWjdANJWVmyGdl0OE6qQVvOc5jMXHaMYGKyMojHLB7WRSqq7NOMH3sN5YQKC3MkxKbqF3+HsDyL
i2lnc0wpPoVlmMlrSprzVO6yQEje/RtVe1Bodp2g3qzUzmZ5PVxZzehjGBybMa0N4BUabFUN7LpT
Ndviy58rSPe+wQ9ZrKuy09lCGnZ2DYB4ndtxEtmRBWkVzaSU0+N++KzjjybkgyteauLoyfCnlCyI
7iw6pADb7C4JJpuF3ne2iQHoRxkqdTZZQhmdwvQFA7Cv4DScNHYgbmjeXmpPsFQgzIuUsTundbH8
vH/2ZbQ994Oc00weoyQAXDpd9PxQnAW7N2wrWrVJdMo5xAyBtr52yp2Sq5pyO5t+Drx6wyvGDfsK
abVvlnGEpnMhJWayqzabN0EIyjVqGgsTxZMSUcybgdFw59iyFTY5cwCdiQ8EoDyB/TwpNA6dHe1E
L3L7VD82lg3rO4At8pnDB1JmnK+ojTDu4XUCzl/x7w3YwkK9svHHF7o3zc/fogp5Ww2JC2ukbgS2
2Y0CWeGmGD7v81lcNZ52acFSDe1juH37F1TQbUyNjAkHsGICmF3EtaKQEGRt2pMIAtyyWYVllKl3
mmxoDAUrqXnZUzOtzz6EkC7FKrFNYRzxxFmuHnXDdi1uiSMoyCo0Xktk4WWeep2Dx4ndcKuQ2841
RHvRnm9vs2Yth3xH8bskFy2A8QrEA0jcBYpnMFYLdE6WnPuz995KQBRMFaEjwzDJEC6o57kO0tKf
MDejhAzLYcR1gdsoIVV6r8z9LUyD0DcjCxIDtl/GUMPfBjhRaovLrt/YIYZmuvUosXprjdOdNQqA
U4Wy0M/HkrditoAvp63rYdgUG8GyApnEUYar8QVbF4GCXaMfX9DMiHqlOqvDiVggBQGv7InAGnNh
lwOdSCfCTCZN+mefaeHkoXDUJ4/BN8didjBVf267LD72v7MvyCE+9/so9l+pTWzNVH9lKF9Csv1b
wC47T3YUpTvD5XsbVD98CAYPMDJVfxuZYlpLlbqYeg+ldk7/yOS9MPSHQMmqHdvaeQu0Pv0053sd
M1FMiVGfebVDbhcNN8UxVjR/H4FH8LP0FHsDN/A9yZmumUL+8mUvogxx1Chcyi+Vyu+s9/lVAF59
12t+qYPC7YqSSLcDKUt2Xa8QosFvTctjQYUt2AkYb7R0F2ZLNAnyK4U6RErFa1ElNOHHQe56yGXG
/iL6XVbHSJc+WQDqqu7ie/IDfvW4LG80y88Qk6sf034cDLA0rPRv3q/yZff065+8Orov0MfrMotU
alQxKmyJMp8qyVPg1SKg8P2kdOGupD2iCgz3UCckOcdlpfP/lThndXngkSC9d3hn6xE7LsCVqcvS
TLeRlzP8XRugNZjFiEusT4WOGpny+EBwI1OnxzV/UxBIFOTfE0Kadop9xwSHrGNYck/Jor0gLWsl
KSQpXH7SX3gdkyM6dIKSur3wSRubqUWfFfsrLBfUMkVf0iezlRqQ0gCYgQCxbn808sczllBUO1Zx
CdpTWufeb/VqxMuwS32I5qCo8inFVEgy00nsGCIMO66asIgiHu4KrV0f4kIymp+iYAT3WVNFLJC+
3FLNCaslwgiWE/j+wkVLngYFFe1FAJNoFOqq4272ZhkX7hICRci418vYlvaevSbmvrcQbR8seTze
lnIUlBf+t8c5TQxSvYXoNMp5W9dbsf1T3kTHU6cur/MyVZEEN7nXY/n9EwDUzwJIfHIqYxXwhxQD
hzI8PoS+mN1DQZ0u2pnKcvKVXTRUhH5IBYw4SwUKqSHlOxE28NKibzAgcjXcaHDEGZKOxYGpfYjC
NjCTvYfMNAqcDzT7iK/Kd/dhBTd/V1HXJMr3iTQOXTJy7Cmu+tV61Of5esm/2mfIxblxpRWBaH32
GDopqy5+/Ndy69bEra1hLvsvumFfcCXiT2CQ64OW479Yr2gNaWbtByFwGanNeBuBM5cyZ+YwdCK1
mao0UmbPpia0mdG4/lotp67ynvO+N+fB5sH7IKirn1/9KsP4m344skT9E2JUXvJQ0kVSRS3QOe7s
gNPgBC44AnTgmCzHtQZWs7i421TQQsJpoO6CiEygIJRkYisW6HZzpLz6b7QSi0OBcLs4XvJwPSG1
LhcLIRrbAawZ/+hQNvw+P1ROhGHYrrY811iM9YyH0wvDpsrCrDVRZlBv/gGUIR9KK5Bc/c11jBwf
1Po9bZrESI35nuOmx4rDnsUefdibUzTzJ7DVkyoPE5efGbcctmDbCxym6a0xxFQCtpCTU0I6sruo
lOlUht5hHvzMK6idZA8oD+rOhbmY7iGTypO5h6n1Sv6D4s4xxjS+qSWlDCDhrY1P3oaEQwoRWFof
hAhUWEpCF4SzWuS/Kej1dF+fe5cr3Ed7b8lF/ebKPoYsWVVeNrwsRHaefMsabOrzm6LdC5EZqxQi
vAc6ElbNOWTtYWSIa8CHswmej4nGxRhH5DPMgjX+8GYZvWjS+rgWxoYFHC4Bi80ZMVCda03PuE/z
wYdy7BWDsFBMFy1BstxSuEllI4V817akqcAKgU4SiCrRuOQvVqlfeEZsW2rpsBRfKlHSe47YOgE3
DSQ2J+wf5BAaza7nZmH75KB+w4YPZ1hnbLn5aSO1ZpD+5fux1ERgK8oTeAfU//EbtRP2ha8R2LKQ
JOMhERPb2KIAhj0grJTe6/Ukn+DgriNd5uSvm5RQ3hsjRbQbTWuxxGBdcAmWjkQ2mbG3hjpRC0az
e4GYLblt6i0L6cgo2Q9ePcvHQYVISi0tYEV724+NRpEqo/cAD2+nfJPKWjQXT++S+9dfB4UikyYY
YVeiAmkt6PdUA7/nQJr52xvOMqNNFkFoILIwk41nSprzmNXut34M4Y7xWtKuX7txZEW4HqJG8Zrq
PdAMBfGNExtpS9y+8txECiB6U985bVP6iINEbaH3f25QDyETBulMoDDbQjG9tja2Fn0ye8htfIh9
ChffAbbAu5BWf32CW8X8dORMBHd1oiRiyDaCM4SGSkffgjrbIfS2SDi4K+WH7ywajbc7Up0BhDaN
V9UR3+v5v7id+7fP1LgvwXYAz2oOLOSxslppnW2cHPZXpg/xPBrPbiGvoAsLPvnNAtjaQ+qdXejk
EAXPUfIzqtfgm7qGooF2DfxH4+omeXpKeHHim+eSWsbhmkBpfjfTYdwtvIPrKMC4Panwi3RrVnIX
q6g4z562DsjTTbaxEEYhUQBmiSLbXvAIDMVuPk3XtyqcIptqQ1XivxAcasyvKlGwfb2bqWPdn3/C
EliVleHzC4c9FmnjwGCrgnZ63XqnP7tMhqPQUiY5jH5reGELcI9quv0jD1lXkzaNaIyYbGeY8Tz1
+ELRciTAKyPRqeJhCGGIwc3qDvpqREiscq1QOZhZH01ZqJWkwj50qzma7Lzk5IcRzlwjx+7IZncx
/Di0E+m5g/hgA0UMg6aoL3mVhrR5r8KD2DKp5O+anLhAhv+yMvnPpQoxU+OLq5aMjSF3rRSI9SAd
UvrI6S511/ev2vDn2YCWEvs/uq/rBrkHJusweXYh6gIrdY43OFX5o7ngzQ+y3UDmaNMkLJiezPxd
qXT4sQqCtDjrXp/mITioomtLooMCymTtYD6F2pER+AxZyBZMoZtFrno6NHQWW4gBPXIYCoOm2uXG
DSYGpvp7dhEQj3M/8yOrijJSYoBRmhtLkd98OEmYuiE0AXJVw0+JegziumXjv3nUcDLlGAOVnarN
EL+YCGIGgy9thf/293sC++zImH9ZQ/61uZ6DKGCumOQi4mnEcGWu0cfO6sQCKx9qvZCSijTFPT3O
P+QTZmR561L9od1t73YG+1zUBoJURyHv5IQ/J57hAhtzM7PVops+N5/60QYjlnKXbBgMgWRF3OtL
LrOPpu3byJbv3xfOy07KTc1V/OGWNqKuDXabjxJm829gp+o8o8MWxRfUNsvvG73qZKiC/ch+PVQU
EYbd5NsOkVA1TMWvS0piE6lMwKODyLbf8ruLIPkYuhw3ilmYGwiEbI5pvA6gZ/on21VatiDG3lzM
xhWsmW14RsvrzI/qPTgb+rhl8rN7iMu9Y08nrFRgPd0tBESPoT2cqxqSCW9IqwBIuPg2pEv3mEFj
5cbEGjzNR5gIWIyKns1MMkiRwFmKZggJu4FjOjeMGxrmCnT651ZcnpXqkmDJPpChzrMWXJQPt+Kh
2ne0GjCzf78gH7bOMSBKbwZC19cIb2pc/nYH1gPigYcvoXIF0FkWCNOqf8+woo/7PJUlI34IYwvk
B8ZK93E41KlmsJw6UnDITvNBqZ177ZOkPg5GTKGnr94ZqBx2IL21m9jwvUp5WQQkVSFBHS1YG6G5
MGzIf55ZcTUOSyH4j+xrDTWyRFpQemtxkf0iPhL53SXk6NuKtQgvmEKc5vexCRMOCB8QAS2aCHen
//G9/tbt+aJA6wKV/g0cTDzt8ik4Evpr7kessz9IcIo4aIbyTqt9E21wiHnhcXbEqK7FATW53ngY
b0dFucDSx098KctDEvYO8KEazOqhugFNx0uvEQUGCIzIh4faVSgEWnuNCZbZMIqaK1xz+UVu3EAl
7MG7HKQWLwr1KZjDq9jfZtpnIJOU5KfERMWo60C9aIhY6k4/lulFPRM9+W6geVxrzjs/Uygmu1bF
BIOJT+bMKj0fUrYM8Yluso43QMMVMc2lTjwlSWApPlI0CnyKiAESYKavbPyqj66lRxZuGmClTiwa
IHq5/AsCFTEphXf2/IgDEF7FbRt98STlQttLH6+asUrIvXPMhOQN1s7oDnwd/MG0sDHOOddDFhhW
7IsWOhwF7rBhgBgAjQomXXvBfgKdwXzOhjfOram37zEssEVJKOlsZuS8Z+NQlNrDkjaFkp3quGII
8gljRQ2Uag46j/39npINUEoJkyv1U2hrXJ4GoXwtrVtUA0CZuh5Ed0O8TkeHVP58UHZlvIHy7y3y
ztQ2lwsq4Csu+DWpNS2sTM2Dqba/cBasIzWeT5cNs5ujpLpUs07qggEjz3F2ZXTS9MUwzLE31eK7
O88QTpLDdmshBK8YJzbSqCqWmCJt1Wx0vsY2Q5ehEistY2Vy/AOWBX5oha+ffOJXeqAgJf8tBvRw
uGZKH+YVFvg1Fx4zOYO9crWbEE4IInxiufaPZ4MyEW5ZxQX9K/9opIKzkO+SR2H90P5xMrJ1XBZQ
Th7zO4NLqfACXpDVi4/aeUpVbXf3NRkmUGjB8wX5mqMn5Sl3Wb06MG9ikCWijeFDl7034aMqvpCf
AT6kUYD3s8QaLJamNNw4kfPM5Py5eNhVA1Ake6YokmhFHfp2gqy9cp0qVN3KQOc7tQNjNg3A7/CG
8vhfR8LoJZt6DVN/KHy2L4qelTH8Z+FKGIGj0U+FsbGNwIDU3EAxaCx3LWiyTO1DjC2nvU3NnSL/
JpghLIWB6v9JW733/L9KzxcQmDQtxNKSikaw/smbdHC/AqIHiUmShkpt5CePyjC2totHa8DdxEFE
YaHtvYJOk2Cgg5aKVi3YCwIbDlTV8g3dGChD6prpa+vIqEwED5Q6tuFcb8jZslNaHSsiDk8XiUwD
ly1J34hPxLv8XUioZiX0D/+z8OnPrcoFIxhicmTqElmdSD5Gk2omJSDKUzpCGARTpjXiwUlQDZnk
N34H66R9SGlg2ogqWe5W4DKu87xB0MethELyqPMkW85n8SG7HSTbdZE9UcZNiBb0PmTXl1FkQlc7
txjrVuXQvK+706EtVJGHqvzwO5NzUsfHZsUlICo87ILz6uJpeei1sMVERdocsWerBF67dGmSZeIG
58dkka2OBQl20UrhGPivNMddV2Vx16CiFjbNSUhF7hhb3PgxXQ21rziI2NsBJwOcr0G4pDl59iMz
E/3YQMXEb+UyvKHLgAnK80PJcA2+hylFN/9xVTZ+y0xtgv2SfFFaDJLUmh8OZOtqCw0TvLy578pi
TFSowWz+6BMRld9oLw/YXOKPah33d4IcfSf93hPmMsKozdzlNpHVt2lvLB/1+2xYZNDOgg3IbWPm
X51qi0QDmBJAcnNJxmM1FfVttjg2zh9mCQf2B9jfgCGCYNTsTm1s4M4e3zWHvUYqOeICKyrrMdBN
ILnDzvGg0q2SJjBktJgAbOOIi5KUP0IMYV84pJFTLPuJ9cKYP54Ktn3ntz73Aa/OCOHuY/v2ECEB
ojCtoGFVTGAuH+Dz9HdP8BWLHM5HWulAhSFP5oAJx+p/ffvq482nL7wjupkXOOPRRidXRNGbyiib
tNMOfum9n6Zx8FQ5vcBFCTaLKBucmoaqG+xebqv1Q3u+oDAJkk5jeqCzgENJCtufZdqv7/phqweS
e8dFxGJhSPyGVwtQw11OY38dThintUS8TuDO1nAA6GhI/e06pYjnLHClX8TxoHTT5IArGoLa9Exg
oQmFVwZZcdMXzmk9CkSA8IHlHB3wBOHA2Cn3II0ITHlHP1LJxe/uaGJURgP6zTSgb5zJBuD8uMPT
uXUyRALdiLMTiVNOjOdyCNHdKuhHOiTUuYwFBvtGi2JjqBAn+sESq5GHNV1LRAP3ClHGz31FMaSA
vpwpE3EhzqKLgNyJFd0fc0J607fglRhnSwB5iRTPNNVxRTwrtdeNjjxzZLfyoXGoU9z5GoJQetsp
cPBWNaoyEBXC7CrCN/FJTYG+s0dMlsMGn5HgzaaV0+Yi5y8RdYwH7oWEsm/LA7WrI7vIDMxYV8jL
WAwHbHB9o60hEYb3NYr3eqwIycskXpsLuzyomC8CDPye7+SLERkX4nyfOK1/w/dOnhWtSJAkgiW/
sJxlZW8hyC2NHkzOMOMQFUX5F1+uchPDkFbsWpfBgok1Mx764rSIpeIX9u61yKPxJNWY40bl4/0m
uyusuDEhM5NdvvlVhDVQz4VTiUFS5I3LhSwd8tILgCaKhA1POPM297Fjd2eoLaP/UxqNp/HaYfri
lZtmTUMiXSxqiqobS9gqaZ9LDYi8IdYp8mmZBCIySrsQ5RuWK0cFgCNM7oR1T5wUs1mkgdnJJeH+
fwjAvaC0qWCOLCgdha9xjUe0AVtWai7YItHUYxOT3ZXxvlr5T1EVV5VIkrm5YvJlbAkdGmkgIW3v
m0SrDb2ksUx6UwEsFazw9ezViX6W8DVwGU2gBDPolajnU06HfYGkg8+Jm1HSb1/84RBSqFBKHS1a
0d3Hkr3dVmRUwpmD66aCalYSD9eFm5PGuUh0Xe7lB6FmVkLaWIsWwUkBACHKQW0VAllan9//DmNH
7GnifD2e0+xsT0Eb5ArYuWqaEfHrxK0rZIssEyPsK0YIxKGWl3Q5wfBpi1VttiO1LGIxHLJAY33A
u/lkB2Hn04wrcAjrtGHREpreq+sWAK4jhxg0BMo63pgV+64u/4An5ben4GV4PCOB09/sLfF38823
TzPylaYmn3cdcUHRdG/e2JeNMdCBYJUdizcPOl2mK29wHYKu6tsuOyu5Sg9MdBoSkl1QGre2sF6d
Kha0ADmXyPCTfpAGNi+1HLtYgTfOPGurYLKpkn2/e5j0Cg7hmTcoaRqBtmXwI0okFXYepJu0g6Pw
SAjTJybtimaB8JgUp7CGXV8KNbe4cZfdfugNamj8bL4uaI6FyqN5yzQT2nrOjflomxuWggrWnpVq
SKZz1Jg4Pk3lsLdJFpdC5RTzOJZOkPlzt1fLYMYVioifAlrR5j1pmTFmUiCte9g0Dk2GWmEbYc5z
QRSEJprNNJ29fro10dy0GSzfDo+g7tnckN2oW9BIvXPhJGWxCFSTimuq/yvgtSPBsncceOk1K6i6
On1cQ0a4Wtu0lj+ua5FfblHxvnE68Ts8dR7VCJcENr49VKPv8oXHI4l3fy2pYL5K+heTI2wKgWFP
SLYBgNUvKdDsBGVOFc6yRGwuDo+eRm53j9PevI/4KERyZ4Zx2gigOf5WsyxuM1QxcFw47Tb9kFqk
B8gHzxIGwKvY8R33DpxHN45izTDng9SnPo/BBzHwwfnAtPnP39Lk8dw+BotmZ/0yjv4rdXU3LTyd
XJsI/c6V/Y5JFbRsspRirrz63mNQ08/JMI5d1EqnR7HECdHnYzMGQJSm6IELaQ5k4oeqHy36kjsL
a6tM76tofaNKw1qsuU4fph9JnguMJ8C8hs3IIB6YMRQXy5aV3Vah9kGRihTS1dWgsXgfWmwh7eRx
UDcgt7ji0WjEe4Su6TounlCP57aL3SeDPIw2ar1F2nq7kV6WyZPugTQdc5ftRonA/RuzPfZO9TKV
TLiymKyJ//xGuA9RB2iqOPjNbQWTI0zoM62MzcW1/9NBqA7oNTBM0NspapIe/qc4k4pkcA4klvzQ
m3CO2K1Rwlv/A8vcYYiGSMuXA3SDaOG6pw8gRwR/VG86y9Qtr/tkIf6tSjTGW8lOZ1QBFX1SqTJN
COdNJ24yVh8b1KN77GCVymE4YQR/0AmyrE0uTeICuUni3NzyQhzeyCtGB45nZdR7jt1YifOVh4ua
E6RlRqbWnahK7yrlVUkmJvjAkqh8+HwK9ub1Sem2U443YG9AjuuH8ujumF28k0T1HUHwrkJxHse8
9l60qU9QCztqenH0/WTjjErjKdvNoxO1udTMjapLezibU/v5mYMmRH1kZ3kqXbywcNO9EgFfNigi
RC5XU0RsxKEvAoLcySFcp3QyIrf5X2szuyNYXWYkssR2ghm6PTkYQYSZb+Ul+QSvtx1SjnA8IrYs
M3wDI5isaXrhSnZk9roydOo3PtGjhH/T7tQa3zyba0oUeo8HNpfphsJ8fdFvqb/2Gn4ZmODzLbun
ls0HlOSp+KnIRJ5XohU7pbAUvTMJwqD4YqffgAlRpeFAA6olldjrX6eOLbI4lYFtLkpBD/j2LjLU
5QP2GK6cUj541ls15ROYp+DmIYBkVUmTxiwpXkZAmOzzmrg7nyV+CHWObVsVVRRFAThaYr2lP52g
5YIH2gKw2k09z/7HNjhHV9n0QGbHdBtzobqsJDyQbsC/KEQCkEM3yyexJDsggMdONQXRzgA1PVeZ
vdS+AiBFBwEdgaNHGGU88kyVWcmrRDb6EAP4767z3iYALy23tNzCKi75T1fMoGYEAuezwlwcz6G3
N2/Pmfkzsml7reVExC1jiLwD156rYq8Co+fNDs+/rJBAeE0IJnpB4I3XzcsgTcgMUhPmsJbaFFGn
anob+bD0SnKxeVzErgFO8VZeFqAkBD5Fx0+46jGo8819BHDvQl9VUQ1eOmrxtIm/i+qRl37b6bJM
rnP2NLhkBPxM9qQ384KbL23j4ceuRL+aGzN79MVDOcVHxmzqcpzSDnOyQ09JBQblf1OohAa3ZOeH
2rkXJfcIZjzTRHIDNfAsd3VlTB9Zkvo9DbFFRrRhvHAdXLVbXWUvDikndw9sH0IQZYS1FOkAnnfS
nlm5nUw6gFxuCK8D0FYG7c/QjEYr4Z4m4/puSOIQIAHsgmxQH3ohPKo/fTcYtYUaDDYf9wqkb4lq
cMssdhof6S5QAq81qgn1/hTWT9ADe1g6VsSMSy000TWTt134+/hSYRPiRkN0ptUo0TbTk7m254xB
EOdMwwyHPeRL+i2feGt39bPIJr8rmtyNII6ZxfzIXxUzo3rop/cKniMQqRv6RuxfxyhwTYlu0ziX
C8ZPUGZ1+CkC2b/syF+iyQ3K18kpN/pjoH88n2m7oVKgefp0Y4I8mlEFPYezz6nGvokUlIkSebEx
4x/kIqc1D3r7Hvnk78qoy4wQcwQJxcYG/L8DDru111P6+lb773II9rXHWRV2YX0rwO3Ia47Tu/lE
Zu7SlpF2djlqKg3QpVpWocmhRdc+AobLPb72Pp8nLx+n42vXBsADEO5wBd9leXSJxdo2NuxgyFbx
AVSmMDDkOjjA2iJDk2RZw5sVDmmp7bSRcmnMTk3GJsiBwuF6Ak1rj14fYz/VqJIeOztmkwj4A81S
Xk/n57qblBsGsY15yxrW6pJVvbg9iVKf1WIZGtJD9R7zQw9lwBwKLBwarPgxWkECC6jS0N2fjRxt
0Jc41qp2LKgy5lk3mSeczJ4QYebnd5WOYYLr0RJ3VexvVgkHA6AW68Mk+NhBdgnxRpt3fD6q4VBU
O7dzWXyNeG0VTtphQS9t2HR8btaXiFF6S9IZe8GylgP8NZXTZH9nEmveyJ20tZ9dVXGAe/2+wUQl
KX0AB5CQUkuOL8pMvWVe+iCfU0A2yaZ5BhK2wtGLmJh08DM6EnHUevGSuHF1783WkAgV13WooaTt
dY4QhHag5dZxFHNMCiHUz10kZoH/Ims/LHR0+qB7RCTJALdwr31u5b59virvERCvVixYMONXaiHM
h4kKCEg9hN0dGRYClaqLnagdV0t0/YIrYWCIyro/v+SuzyT3/GeSrcmrMzxAtt7XVhBSqQlMu5of
D+6IAtCij/Xjo29eZPEAFOKmI00pyH5v3GnI1PEPcITamJ1zGfxKZNlIjbg0KfjGWXZHowFAyNL3
FSO1Sbu2WI3IcMsXpLvYkuwWFu7gBOdJWLKxhSzbvA/8rB0ZlC9A08N6OOZ9GmZsJf11WGPOfi8Q
oCv64e0lROzYbAcmd4XB6sXx9Vgql9PhAFHOOJhxu6NueUhaoawBkjRsdLYqtNHkLvQXcHLYjNOy
w4bzZO0JKpgBEY95xZqkOMoYXlePRLr2fkqTWUFZpWwrSgrfoT/s/JLJSaOR0tiRzbX/3q1tTQeG
UW8HRVcHVLtgwX2Z20dfchSYSLA9L7C7YuZV7q7s3M1eEvqxm/Kl4hyBANPlo6kmRaam/BKUfGMm
d2NZfn4Qu0jdO/UAJqnh0WkHSuX0rxVQmwyUWofBp9OdOBX/DSbqlStdX6d9slGiGMjKaSqd0JeL
K/bfDEkRjkqCSKrNnXVtJUAvSF4UdBVNvmfsEUWQHAke5heUq9Yfg7bKoOQ/ErCh8EVr67EgAfvJ
a15L7rQOm9MFh8rnlJLeVV7dskKOUyzQ3JIIZxdqHkQJTLybOLirEmwGJ7ZSG0gRc+qGoJ5dc4La
NEMrRRFhWp2T5s9Gq5wPmVxpn7t8lY2lDkYFIQfVlq0JjzCrFyM1p93jjWbJP2QML6WlAnP1Fu6j
ZmANes6qe/qraa5tkn6uHfl/uvLm0ACiB+Ft58JDtcqKRREs/fgcGqhtUiOJtu7vOqT4dTVmkY75
kINhxm8UheXy6nvqz/qiSlBsIHs7IxUwYNy7XP4UeyT1bktMzw4aPcszytPxCckS9rGkSNdD+cDY
uyohWjRHMDc3qQMtJbZCoQCyw0ml7oAguWKbakzVcIDdpVRCvhA2/c/RZbSfsMS5ofFKiVv3MGaV
w2N5DiuHkrQD333kUJclGfGnZ4xtAbQC9Nji3+Zl056WQi4LIyVqHkX7YAuVV16SudjiSeNgY97o
SNh79NPKC/UPQE325jd+zyUgZjEyci+MH8HvDPrTJHaFIn8yLKvVeed3TS57hqiAqxrK/PsedwaY
0Tg4Go9beTY64n6GTTSUS+Ncp7VKyb46tSm4AEy5Lwff+eBFCHtK9y4T0DGoI15fmD9eTEiNGlzr
9ezpZzu3KelhLaQPbfZlHlaDbPk4PYOqFKVJbqp6P4sX9eBlwIDF1QMF3760IJYLsvfeJ04lr1gh
dfTi7OHV7Kknr4W1aoLhbuAaRwjKnbcQOfSa08Ekta1xUxn9daXbu7kwwRzO17o8gRdUd9o5bqV+
/lfa6e1IaKK/QU3aw5Bc9wE04vo9dKC1oEMYf3SScz/vD9DLl33pDfFHOr+cPVKA75kXGDylLrKS
gZ0r0Cn8uAIyVo7CXjB/1idX8f15YzHs3JSmx4YdDLcN5lU6Z8yNMS2FYfzYbFp+c1TDb69CpAe+
SYO3TBo95bDQpTNNQmABYiAQb482mveZbTIzaxuphOHUquWzn0ekH04knd5ZUc8SOe6QiYvvDqUb
f3r2TF1LtZNHeExIYNo0U/cRthRUcHqDBHZT8FAA1TeOdhM8d/gLjR+vzeodCFCsdh4pXlFX/7gR
rTbOgr03pKk4KW3W3oVfaoyS0dtaV9j6BOAHQT8iGtEwi7muxpo2Jai69DzTjhroN3TKseekf/N3
sziCPowqrFNN4RFfD02tf0K0gf9ZieNSG5E/ZD9t24YKuq04x6w9NAkSqTtKFEjyshnZGgv9spto
Bhu8eEI0s8VMtT0S3OaAxgYgyeNGkhu3OYx9Xyfm5nda32VWhvTIWISjql5gILmND6dpFm2untGd
zuOSbpIsFa/r53zCxBt7+xi+wYmwQ50fSSaajVzX/qPGT/olBoF5J4GZiipORb0IHNPJ+CaLh8nQ
qGqAkcIScgQK4dYcPd2xKaWgFAdgu9FYNIqbwetGA99/Vq5zIH2Hh8NNzlXIbCVFDOiuz+G1nEkB
WyjFIfFgijV2TjxX1fMW5+7MQA6HT+y1kuQ/mZedw9bUxFJXovpghy6qG6cpiT++8KOBIvyQSJca
hFVi+GDVsjPuWq7qcdEah7r3isdbZVn8ziloGKTAFrMjMLUr821zoBZJFAWXkAJ3ic6qhyuAAyXl
7TNXHzrAh2MbrTOY9yu6sXBmiyXlU5+3m/a7FREJzxUP/kHkGMNQN6UyCPa/aI+E7VlOweClPHdW
IshYfkhgacVcjvKnfZt5weUcZlnURbgZp3TAw2piZdtKN/dvF0k26qQ4DM6zNZgWlBVPaDbVR0Pe
t6vfONeYOWSpF1QBa/Y5y5G2n7uHuI4J37KVLI2TA+F+bz2K+u3vVXRfyCjhqzxOvReYDaLcsQhp
50+exGD5WovdnZpEbpkHCl8/angb+7LJYbWD8qkJLu8+WMFehfoQlH3YkUFHw7TP6al+zhkp+Ij+
ZiFr7YkmbsP5tkqlmSGDKzlhWHeeme78kv9Uf6LXlCycICbaWRHulv7HjSD5cgtCdXVI//nxujRk
3z2YDRbAgp3JHPzBnys4hcO2nD9hRq5aa2ooKlRmzl/Xe2SoTylAbzqrIk1vF2rCYNg52AafeLui
KgcIeNRGaDhOGIdl2JSiFxiHhzrWhr/S/7Wlm+iaZk9SQS4gDgeKr+IUk13Fd226eKEWext4bqul
IETBpUglipAbXy7ceCI+CHEv6fVGrH53/45Sqtv8Ss4IbR0vr/E4oDEFfVJlCN7FTUMoPPxBJrjs
wfv/idUXFDGxjaLGYf8oesonBSt4fjeyt5JE46AME1XHOQGZKvGiHjI3zmdDQtT+zuy6QVFqHTMX
VvKxgEbto42mcPY12WMkre2U0PpaQsml0zyQERN917HqPnr5izYqPvPFrm4XuLrQC5IrniuBRchw
4kvqjSjMbDyFbxwkIiEnhVa1eA6AkXYCBM9DpM7lecq2S7AgW/OVRgiI0+8nq78wDAwjV2yrBtNb
gHVmeO67kxukikffXiDlQtEJGcQwd1JoE1LlaFg7w9IRIzpCL8mONlxH/dn3I7yYOS7qYKYZqBsI
ZxDWNXjZ/KeeP3ndTNF1RgMT59roebS5Cg4N7Gj0sGrvjHbY0kORIhBP1GIdPaS69q9+n3mhuSxK
76iXUNo4BiVMJvxPMZpb8/PkSocF/cmRuX6Tx5HtukuAk5S5WBrENOuJr4x0/F5TDpO93643prJM
O6bwFg7QbpgTHmwPqG8LYqi6ny9VRBsom/N9yPHVoypxdRyRL4xVnhppIqWMDMzPy1fooSiGRnyj
sp3isNoWuKJIHGuYssCEQXFHwYPur9YpaJxTlbsXZzeOcg8lAR1FHHTlzgqYNbE5q3+GdYyBepdV
hk/BbEzmwBGH10+rxvw/IvqL/HfUVY+x4IMr9PdjZfQWmYXY4xacqftzyfnN4QDazUzWQcvmfkBO
jcu3YvT0ppg+qazJP1Dj7H//DJs37yCRFnYE5OzbXc1GR508VHywREExBIgDkrH7hqXrGlxFxj5t
hgk7KjKXqxUFqVIJXSgl9BzfkvlbfYWceGPU2DVDkMpX3P01Vzx0OQaTnBnVZrs/ASY+mts8tF9B
rEad6/eY6Dyxtecv9qMdxK2SWA/pDl7WnRx11AWy7PH7KMUiYPG0N/bFlZ0oxzAYeir+rv238uX/
G0f2HI79xQBOupf7EqONraijT+DOFZVWrUEHefszaBc5xSVf2cYIN3pDymbjBEdViCAe2IihLpcP
fgCRB+EuJ4P/QJaE1okD1jBbOXBmXZ844U6jHk2ZofeCInI+XtB9+NlTSpjUIc99U4LZjK5FzDa4
iw/+teORvVb2MJL4uIg4sa0ezjpzlWc8w5uhZvc6D8fDB72WuQW+FPm4COStm2Fbcem3tad/Wjau
QxvYUwA8ebmjd76/VefOIx22jtWS6Xq7xpa/yNioMvriB5/hIXUuzuxot2Vd20QzwR9dvLheTXy0
SMKQQ7z5lu3lMt/rPgGkeryvIs4Se/WDQXReF70HozhYFWUHowkqHIBdOX7tGb1nlyzbQcGFXquc
5GjWFEk+k9w59kkYt5KU0jAk6TSybpF1xmLxWMolJN/2vkh8ESCKnNpfuCu3+es3zYtnnZMbl1hl
MlzpAImqsO9YHhP1o/MV5+k95NirR18dkY6S3EgXoiB5rAA3Za92M98DgebOtwcHzBoRqzir8GWC
hZGPf6uw0PXx7m18jvbk0oE4nt/xPCcb9Nq/f3pbdTcQqn1jOvdPpjIh0IwF3IY91GqiFUEIrYgn
STTb5WoIbgsi9/fjjwD6dIGaM1HiTwpBarxWENLJCbk0rmk2Z4AtkL5xpmxecmgMvJA5mGx6qEWr
RzSEGjttwgbIXogZxvMdf7o8d53MzDaKxVHThi4uYHOowz8gXpCZ5LaG3vzti7enwBRiZPsgE6fA
klhG4luX/1HbALov+kFjyRuPpYqN9B2r3dj+7h14jxDABHHqQA6My3AvEnWeTMmqL/TXjY2HsafO
VxaVIsBQMxMindZmszxslYu1i8RBlqKD5rBdU91Oo481qGLfoblW20bjZTscDmHmEyFj2cp+tWlh
/ztODJmxT09+aIbdl0RIXb2LeKib3aoFar17YHQ36fzoRlZaaUdKyQpCsADm5DgedHUtaGo61nTi
gUOBIhxmsmjBeD4shS/3DDC1aaHwEOrfy+lSkfuZtahVQjnj79KTp8QS81iOyAJ+OW/Eya0CW0DP
5TPfwgr3Sz/9yy8JnErSa3H58VBruUT5d6a04j6W1KFjVjfojzcEY/ZGxQl6lpJzpYpldlwbVW+/
CcHrp93jQE4NqcKfhYAu/DSgTi2O1FHWnMCEFXZ0PWzdkm9MtlyMpqS9W1l3c4IB7eZzjDVNa/7m
u64AlDcVdZFkEj/FDkCnGXblQlNVm3oE8ikpmVrjJhn4sT08RjatA/Estz7ho0BCXkZkj3gkKrHI
BX8hlrw6ZxMZSZT4TT7uFJiZlTIelBry+f+kAvnFfDpL8agWwSALI8wjo+c/d1xW4kP/Eb65GAS+
FMN6HY1CTPJ35YhUpUqI3dTjyrXG3Wd41NFvJr8dDmmINGBZlKsQrvivhD5H3Zs2DLqKm3/zUw6K
RMsShXeozAfoHDuCx793wKlbGCQ0XnwoJQSkn8Py6tlU4X8YhVOCj+Izrt42uvCOcoWIOykd8xqJ
vsn7L8UNr7RntnV84pTIsFU65zJj1ukVEz3eyptROv7xWSpO9SsjCe9Rzw1cS5eDZE2ONQO+2W5Q
9KxKFlZeqLX4xJ+ix7b2GdZgL84GtEVi/OdEBTlZSAs5UDr0HeuQEFIFM8B0HLyFhGKcHe7uZX5a
yTak2XSxcrGYPRdAj5lbuqDGAamYDJwAylNxFzWkhd3st5jOmn7MTxG5vo5MRP/IWyalV3kM0rw0
jL9z8X4ulMooKaRKx4868f+OsCWvAMWlmPkQSr0WxjFqsVq3GMsnBlOQLFXnXZoadps4AxpCut31
h7M/h2qN/jLgdmV9Pj4RRi7ZORQ6BdJKsWZskSIxbCCz3E5VSUdx82zLw0qAe1uRcA8rlGudNrLR
hrEk2h5rpQAKtYFHDN4IXIjyR9a/kiOMVi5xYFvF7XsxwGcVXwhIlqKMMJBbVhGweaGDEqBiZaNi
tK3mupkoAs7AemyavvUQ/dMsnG5+kfZLC4XYvzpFI70hWOOe5OoMxdJqwSTR76qVXK4ErpR2mYKe
fo24fSBTQPYx6BSn+nGpixxoxdwq9lqm33m4LLi2f4gHrYHJcSnbeFD/2MZShNfGoK1SNSrDs/Me
6NA13ys6HBzWYiXCRuJbGEHabohK1UNjGaQ2rJlPcm50O2CTQfvbAJDabKyjCk5RGhHLpqbjUOHS
8y/sgadZFh+8RhMw2O6xsqkGoq2D8p6NXGVJXQGkwZ7S8KgrnGWmema8WVmibKOYsrLLTYvTNrFF
qYptxO2PDNMJeE/m9yO/oF3nhwUvZctGFxMFJIWjnIlhY7DNnuteVdjJ5P/N1o5zrzd5XYOsCHv7
pJE4SVbNL4byrYw363mZhJXNLgKKmUJKJsaA7FhGfAUaQCoRXBCcRSPJthS/Cd6XKO4B0gYq3hbA
JLeWe1vDRxAWAmaBPb4Q1qH42+BbvAaBGP2FDwGUOfr6kMA/FdtWfqCIneicoUm52JizwwvHgf8Z
UNCk56W6SDzZZReCr8UKx4XMQIn4T5kOAtp+WRrIJtiaXr2T8v7cyLMPmFJVodA47lEER4QcGMa5
VXt80ptT/+CNWYH4CWCf9GFfooOPV0ap/LUVeSvlh/NdNeVAai/GqNsJJ7/RAC91YmHJFFrD4M68
xaVR2qdhfBp+Vi97uouwHjPyEOAjObuQPIwGWN0V54AHHjrvQcIQ4sShtUO+w5bV1YLrZs96dOjs
I/08SW8iRpD24Ft7ez5Km8e+9msTlDFhFNTicdbUYvb7Xu2hXvJ6LhM0iVJR/mRzp3AQDfkKMwrT
W8CWZ3k+JeDkvWUpFiKX2OVLESzMTzGRfT4UACJ6r5gG6bXjWmqXH1qkhk3zYRGEo0AEQCgKOjwN
/xqYCRypdtQ+4WntQi7ih3ZHuZD3R7UvE3AQzigHLeEuaA11d0MXiRbFZNcPOj8wWDEGlBkC2Muo
579tuhM9+ad6K5La/vUSr5vTGn7e2a8CKh1bqzoQR91601ijVrRiiKTTafDUAFBlf/YZRK6rXDKo
YoxnWvARpbnSRyR3MmXZmFs5wvAGY9ag2RzkbO7ff9Vf+bJLFcWy/fM+s4wdEyTyrSyKijaDiGve
uzV2sWFvb5GlE2VYxA0FrE9yl39U22sD4Z3ckcbWAXpSkspVw/a8ILblnI15wYrf+Mz3ShQXqJmA
/tTSxq3sRYkRBkktnvUyJ55oDL0v+Cet4UUotd1tHlaPsrAZHrRo7GcR8YAPDWl6BDJbu2cJXGtr
ALWQFydWG7iJaO8K5dUfnLxTIEYbayMp+sfXsW6qmgmKenPm8d3FM22v570bLuwfOMJ6Zr3i6Ldq
sc4DWH7oSWzYb48FF/3YP1FAMWqYONtOQK5qd22pbFYCR9HlCuN6h7bZAwa7Va2UTnRZpVWGXwMI
6Rmb0aaeWQawyFqpch2gMeOn2kNVsDWDnTOUciVcQYMbEf1cWzvvIBxkUFgmSYg+m2Ufppm5gtce
QJvtusdaaHesOi2nI4aewkgPQ7CXVSwbJlTrI+T+NLC5bd+crvuc/RgyYzd3dyFEOuU3qE3Pd6uU
axtzXQ4SIHPtA2GFu254OuyV9EPaAoyytXlgTfRbL+chMBHB5ChRoeSZ3ALkHQvvXBsBnqnAELQB
kisNxgMAuUazTAYHdRfYmbfFLOcctrtGYCv16ffQaHKkayOpgX0W1/J3utSlkTenluXiF9bK308k
hWljSnqKyhFBaj4LdY/OGiclZwHCa2bJRJGxrJcbuMoeQ2IEXD1YVVd6kgElULGoxpL1ScXRcA2P
5UEdFIvPZmutxPMoT9FBIWsULH8V7LLhSmNemW2x2IS9a++LjWyEr4Wt8VTXtUGgdsskQSgkzSzC
9EbxpAaY1kauDhH+Ns4Sa9SwPUoJ1F9tavLQWzYd2j9LelQI4bRzx1PtvOA26y4uu5pULdeur33s
8Cn0Jr64Cw59DVJT9B/QTGtZoS7MuX4jv9hkbyjTnW0qEMmQjjEBhkgLeGVAkuV4coRzPMO6x0TM
lMq+PPFJ9HVv2xIkfz8qcYo3tw344Be+fgbyHwbjBLBExb0eo0qCLk1zWqa7ul5Xf84FbQpxL6lE
OzgwcU0ieXA8QZC8YCU1Lb5XcDfrblVBar7u6KShB6PjYvp5S37yYRWDVqe71abkYhmUPydaVSKq
kF5upYtSCN6qKKyApSkOJp4weP4jGCDgdvpIUxdBzuuJpqLyuvkcoe44JxIMP/C0ISwqyFfqA+2N
cWlcztwHevcAiprmKzgorvVWfHwUQsFA9O8H2bM5CNwOvBQQDfoeBXPMF8nWejzlWehMB1w3Y2xF
Rimn+01GYHz3h86Q8Y0Hp3dPqmsl1v8enX6QLMqV6vX18S4Ko0YjKRaLt8GPYAGNdu4zqR/o4Q4P
wv9j4Trf+DsX3PIzu/vCHoW5JG1WjK56WeEOr6ESSORJGyoMWj6zukRcotFdTgEdwR1HDZ8qffEv
XdT3viZNISKcxhgCJ+VdO0nnK0JT6pPGCp4wP52SGgv9BSPAJVpIC4WGx2RoDAFayPiI4Gf6diWF
B5mZBY+Vh9aMfootv/E37djzYXSm5YoK1GT/8JFsm991zAyxeJzwh5cCxDjN2lI4o0SI0Gg0E2jf
VVCSzq2CT892MQvR77sNBNMUiVSd4BZyhmFRc34WsAk+69qyo1bVjNwAI34nhx4EKyjjOyLS9E4M
aN8mC6lwkjkjJSwp7ch9fbKGq0sG/AT5kqWtF6K6XveXDa8Qdy3sx896eqOKV2M2Vpbr6k5yjFzC
3eUWkiYAmGZ/naoJ15OAuaoxmGS7L4U42R3v+A4eFe35J9kG2vAz3EewleNsMF5enPSF9XmMaP24
yulBVKdeXNXUR60xVtGPlPsVb05Ry+NE+zEZXjGF6Cmwlv24WzHzYJkiaPPSqINH8lSKxao/qsaP
IVqo5veinT/of0NV0EnwmoFJHm08xDWgbRPHggAogK1vIAwOm+hVuDQhyk66k7L6z5A4SbZHIx0N
7bxEdwtf/vMrMQDeIsIeLoNO2siW9NMBKY9L1mR5mskVYEebWs4KX/hYxbsvBJlI8UbwvnVrnifc
lGFIUo/vgK0DZse1Fsf6GEds121PmbfguA8bRNlEseAkQkXNpkz75G1U6SuScHVkEa0zg8KpALNK
Fn5yhp+GJJSV9ICVlx5QcVXSA2GzhAUriiDok4r9+FiIuf/gaaCFXmwaPWFcNZsuZH+c2hnaOrX1
sP0KgGEiRHQ5n6EmqkAe/Nx8Y4yCrLdzIe8NMhTUI0U4x+EcwdLlqmQhC/JNWTsrYvRT8MjWqRg1
5k0bnBOyTSyHiYBPDRZoDMY+kDNnNFbRYZ2PF612+6ezD9ie+HpP1Dp6dk+2QODvOs9zmTcI0BVz
v4qa3F//ut9gjdahc/EBWbTgty0b9LEmzTHHUVRo6Qpc9J2qRdASJL+zScfHf0t1bYVxyVehDbMK
zG88a4y5fBApGWs9Mv9Gn3lill7/esco+AaQNyVs6/2IVUp6Tp1IMReXT0qAgKsTRIOh+54TXlii
20zaIKRmTVCU0a/zfhJXLZZre9+2aBb5x3CWPs1mnMe1l+9A9H0whTR2Mpbjs0h4fGt7RpX4SNAW
oB60ZgNYpjW3AqsLFTE5gvXXKkOjmhaPUPlYbXKMfsFPjmebRaGKll7kAk3/6+xGO5heA+ihaNng
TB8nSpgQPD16LOxYGcZ2jRWXzngFci4gyBL45XPBLOAGynzKiR14Uix0BzE9Ax/4h+GZ/SATg2b3
sPBlOaxibsVtO0ar3K1HfaJLFXfoR4zOcCdyFuhTKaZLgtYtnPkfac+O8UcCXNAJ9d88ZTA2FQKU
vKCJ9KUv1STJgkVjBjZEJyiBqK7JTgRFaV+V1GC/B3URfIHeoDhs7wIz7DB0uRkhICGjhRjCI3wp
ATwPRoihgTznQgii+wsMCR01fHEuxusQG4J9YxdwYsdB6O3dBsi7o1JJeihJ/6V683GxcY/rVdco
glYvNUe9WmCYca33oIvN2+sZBy5Nm5AT3n4UsKystmmJT49oQRowJsjPQHWKVpkWeS1n3muSO6E4
TxUtTt4rp7jFQ/DtC++bIgm1kdwIJzeYEPsm10Wh0DPwrfEw1MsIpur7BU5/0ruwL3+XwciiLtPM
Vdn9OXuFS8SRPk5VZ/tSfzG7U5kU+LoRWuiYsmhHD21HDEl+SSysZxGP8DQlkwaiYA/O/tI2Yrpe
9hR1BDszkgW+puZzRETPCJfc6RoyCGnD2PaZ9scQw4hYy7OLjW9r1HtyLPdu0MWFhsJaOM4qGwNE
jHS/vybI9Qq78f+QY37VFJNu6KxcL5Qg8PcujVsI+ytSXC23nKvbHkhypLCzDpHOxk5LAPLbZU4j
p7r5P7BdwRnUs+RE4tDqT6QgN1RZphKkshnXBzYf5P2aPaL0WCKDlRLEa+Qm5/8T6Of9+siVKpLG
a40fM808nCMV0jS+TOIvbtUJL7XSTvPnMnaoHu/6Zc83tlTL+7eCZZytqj2dUlcHSFbU2CnlAhU3
baG5Svhwvz2Sy3I6SS5sdhuNZq1wj21DWpYo96ww4ZUYlFCTo397uVf814LWvU3DZPNMrQhkBO5W
aY4LdaCKIfmwuzobIvFBrjRaEiJ2e251AkuSvoH3eXUqhiqPMYR+QjSWXUVNCiIGEOtVVlKpdQ94
IUl/erio4ls8LexVvikYpT7Z7AMXQ66PxUpzLJRJFGaxZ4Kp+879fRnUTtrTUFb/d4bCmzDLT1Pl
kk75mY7e4nJS+3fOQndtIjtFKP3FeDjiyb5LMwwPBgT38CZ3IpFY5H2I2NQda7raxedFB3zrJEit
qcrIwXQejxSZvP5zrfY428dZ1L3+b/Nx/5DqXC84OE3ejq3+DAfstqPUWSNrpS0Db7mYc0SQY1P9
7HYnHvoBAnHJsQHFO/IEIhqKeezaP668KtNqYTuw2YQiKWhnjhg4E/yIcNXCyQqVx5xsOGaSpFwq
HLswEctLd4sbc08pgk6qWoTZ4mfMLIAQA78Ies3vZ0BYAqLlsxl359BSzKKNGGqwMKNvKa3Nyj7n
JRsmIvrlR5gW+cjkNJJXsZ6gQT/6ZEXRPQii6CGYERqeAgI7kVp2WdnPY9xTcajbIOfDD6J9hFEN
6iMb3Zspbx0yxuyKBy9X01CeYUTW6AwNQzvzSsVQS6vlC2ATCeY/DqNx+tcAamgKyUhydlVShCWz
PXcM2GCkvFksRB7gnuhujP9++0hqIDWDDT13znDcacNNjCTVZUPawdmeJipohJQ3RXbLCaVO5QPB
kswxTLzYDzfVsdgZZF+QMP2hJuXq/NOEvoHiu1UbinYOEA/usQqmdopmLaCtW8obKvRj1ob58io6
tuMqShW5kZ0FAXE4d88OZdl3lZdTol5g0gRE+PDLLx77ettoVEoaG/c0kH5WrBR2KxNSdqsqToJj
68pfq+V0cLAfS9q4pX3sELSNRoxx5HE9tZwfzN0/j+QfoTWKodyvoUaP5l0bxWgJquDkhB3DS6xC
U5gcxz7VRSnlSNEocALISrdHc38jalrKXjMEZ5UDQKUszI2QzOClmapZAF6AKIMtIfcp2EOxeqoN
P9CoQdlgQLlQ8VRl/WEvPS0i2IV1mI67B1ZMhF5Qz1+5t6tuMaUm6Y/HRiOVnGwsdSe4VSUl0iOY
6WjMbTWXDYcWU+OQMzopsqJxxNwXkD4h4QiUQW+0wIpB9dxag9lWFu1vP68WCo5fSIH+Kgk/AC8I
VXvXX/YVEhhc26v9bUPYVYXQ/LFcSLmUkhSS6GdFJ2dO1PXtW0W1LNAtL/cNdIPH5c3oq+vhduId
rd2Q9O84lUR/1ukZd9K25N9uKSTTWqvJTF2vD0dnw2xq2+45vEhze6gz4iWBOHyNhiC2YHNnTayx
2BK+KW/Yix2GQ1XQ3kCHAhfuQb0ZRed2EjcoiDtGHMQ8dhnRMarRq3GYMpRkaX9v+M6StCkruv7K
pRHvxX7PkGVpRvS6Zsgab//LmB4kn68SoOigXP52adaVw+/Zc85pdiNkNmwS9C1wzNK/PLB/ykL8
wSD1QJumtJAiTt4z3TcWLQmIcdAWuLESpI+YE6MgLHi7sN0LnUye8u30gkTJukJeH5KVDH2RFb2l
eMUbcOD8YbvJGA39hXJlTAd36C4UMWRYirccUio0uxoD4YyQPSy/sxc2fI2ZCaiL1JDpUU6CCL7n
klJqJKd4Cu70YkcNWrKrGrTjc0TaWaldG6aTQcUIdMPq5W79U5ORzZIzF9SWtCHLefMUSfuWgxYP
4Yg3XcDMP24bSdhCDNU4hqApbmmtL7nv/d8SMcfwUK/bzYXImH1Kt8iaXmuQpcBnk5EzIaMzPDRi
bDcAP3sN6u5NKUyOn9sOKLwRRRJdpqLUvBvqfjnBS7h3Az7Er8jnY0nD4XFeNATaSCf00QivgpRO
CEkIj1zy6MoLAV4/Pv6oocbZWM0MUzVy+4iK6n8B1NqngIxw3AQvoStLlU6JHLNc9jxzc7f/BtB+
tg0S1BcODH8f2MtEc8iNjiiauM1kkZq6aVP3wu+avv6GKF3Zr1xd61PVA05h0Cy3TD4J6ZC6Set4
RwIwP70bfhsiz4FEYUfW343vJP8j5lIlcXELYT3pwvNkmWAE0daKoDYx7CIJOkNkDBp4eTI0LaT0
JRE2I8BdwGqukdHU3k7A4JsslrMnJFfniLAsutzjpmxOdqNYo3c1sjXI+8LuwOHR+EJXVDcj6e86
vnobBqLhweT+QzVIcWj2DL2EQH/btVJF3RWCgS91vI0ZDVUJvDtBjKzzkD2Rsh2Oered5EGNiFrC
KrISscgIKhHF70UGZa5A/hhbqK39u9+gNot1f5JG3mx6Vx6++yfsR7Y3fXSWOLVa5kXRmhWSOc3V
O4/5daMkfKS0Rkehims2jG0r+TWMwd+Yn7F65WCAHJBzu1jXL+vTwgBCUT0SkR9HUa+LaZ9Uca4a
ZoFE47D017wJS25zI5X2BUrZAGYm+gxgMjg1fiCZwVgYX/+13L6xivDwrGODNFkeIfZPrOUC3II7
ZTZbUVwesRc7jTcA6NyGz0FhQoTPFLzgg2tHOd8tvGjy5FQDtLzV8recuU2mDKwI6BIRI1KxwFql
OdxsUtn5pr6mbN1xNZjX0cva1tU1yVwWH4ZomDBpzJ24dJyRN2Ao/V1EinNjM1Eb/EV9t3+FgZvz
TCmTvYFniV2nboFLmmBar+eELKFJJmtA0LAtiDdMSjPhpAD8YP1SspqCC6+gjHV8k/3ADj2Opgoy
WIZd4VYbZgRO3w9fj+biDDg2dKFAPr4WEIr8g5hZJxeCA9Dmj7dxB2/Z4uIkuXhmV/BKhIDzcdLf
sV0RLxF86c4Fz0kosuT6qIdO4evpoCk1xi1LUfK6hBgaN4CGDVeg0jS/5vGdr8fVT29afBxMsP0d
XXKcwnU9EjTcn5+OBwKBgajWdmfrHgpPDtjPiG8Uyl654KpHW8Cu0fw5g7HGfGuxa43oNBJV+BBM
AHngZ5pyJ1YEyNn7bcnJ74PzhIiWx+bb5UCkAqx/IMGXZFu+Glzn2+mc9KsoS3JfHCLT6jqt/wgo
6E9ESmv75xOfk8HaL1Br2vo0Y+wTaVK4oWpBjiPNcwnvnBahC3JWc/M9YvFDlNz2YTQheV39xvfp
DlyGjCcDwgsrvB7eHd+70k5+Udi620jCA2/1WjsZ4ElvZzdYM2J3CR0stoee7c3FSbnTFSJXSfJ8
4NmTZrNZuduB39n+eCzV+2ZqYxt82LBm02Pvq0uC7EsZ6Ngd5mLWgNqqMIClilCJy+EAfTwyWMgu
47oxedBswC05Sn96k2wJpiXGK8h5QyM4W10fMmwddOG7oHJRCWlWmjcv5v5l9Dxv0webTx/DlKYZ
Wz61gdKwyfJsSBL0k9gfp01SiLKsNl/7ZkrIeDT7jpZ9MA7IeG6ag/P8IeE7qIour3v3O7CxXymX
ighVneh06JT+XvXYkpd3hcqB7/LKeDlkWauFTFN8YhT+dBEaGWJNIUGeKJvDs8Sy5t8FGQknxmMO
/ZtBe9psx/2wUBDmrmR45cdIW/IgImquSNquhJgSnU2aV0JvgG+0jHr+WIu/IPfRHLOErmeL8ReK
1CxyqtwU8V5YDPiXua/RDgohkC6FnCmpE7dl2+8fWSBbww2t/A9TR/DHU6ZYq8yHqlTqIbNAKcG9
cc9XanQyHznYraizZR459KLZsViHYz1igE5R8zACyrcu2na2/zonH6EGmxMF2aIfBGGRf3iqUNDu
5zjdUuK/Ed3lLd09hZPLpPTEZL8/1m0onubKMjWHxOCqukx2L+hwg/Cs6dA/0bO9oShU8Id5llat
aql3faBMSTPFX6B71WI2/g8mZsQ5gw6Z0imAHhX5ziU0t/rinY2xqBp0+SVv1BoYcWLoI9YyaMy0
9XGDvn5Oqr9rDmUsKBoK5b+UGC1RvuWwCJQ9tLD7rRnuLJiXLabH/NFOTVzbkk6kHAZJdYVas4fw
ycooa2vzANyEEm/V1jyGDQu66kW3rZ7xynokgz3VGS4+I0Uap/2suo0FFSPptqajYCLSTwg3Hvnv
y04BRrziUI7ByjdZnksGgJtn8tdWMa4PkrykzzS0UppRNVsSOzYqCchVlXmlKaFY4A/viG9hTDIX
3JfY6vfNGM61Sy11DQ2WSEzmjNDCoQItVy23eONvHh/VJ8xstHk+++1eai0GSbt9OH2K0icgfZap
hTN57O1Ns7lP8xGEzvPpgdtXeemRDnKvHwJ9TZxKT2EIRfevxzJbKbYeP/cPyxgITuV4qrM+BSpA
8RkKL4wuuecDsPOamBuqopqhfvSTanhashQlK76LVFfVqxA/cft0WdD+wko/8/RHK2Pij8UObiXb
ebRKBY7dkrT4g7GRbYzIkCJ/ILf0NBYxGBoInLK8B1y4HFhvGzvAtCOWbgpYyASOB6dFP/z1pr2W
8llO1wUYasuoviu6IaPtvIYKr7U4Dh56eZ7tny5UE1Z+L64yaZXnHYcn3bZjvE2ytyqsDDcJ1x0W
O6+Z/4lPkpWs9Z+KTKxN9S6wB4s1+XQvpQDVLymVdUk+J5TSHQSO1vgMrrj6upiELa4OuEjfNtSf
JO6om3k1M9g4qffOjrmZ0jpqaYuN54PG1wjr4pw71H4lSG3cmCbTctdIG0Hlz17U9iFaCrfklex2
zTu1LsmrarSHl1fQ1m9nBO2ipkN4YHjt6BIoNHqCN75uAAJFz64QcA/Y4eyDWqzMqkhRbf0zeZyG
d3ERcFrEHaBNguMZsHbxTWgDuPbgvqJqSSVwXR61qZ+4gaz++2+0T8QQgJGzJ7TQR5Hc4T8xvFme
q97jbWTEV8bFmKTiaPh3o9BcxkztRvk3x6fsFUpIg/EhWk6kWKE+awPgGTLOS7Sr8ctQgl/vjWPV
C+GhreZd694nSpin96Pwmgzpl30a8xQ+QlrzxyJqRzW+Y2rYo1HY60urQ+/5f65kYcSieRcYQP6c
kDT/FmRwDQIZp9stv0U2ZiPx+dRlhr7kWwUyvv/g3jWreGgXtZDxxLRyxlKsJwg7kBGodQg8Wz8Z
+6Jy3NHy6FwQAe067NKwM32tfJQaX6TlPpg3nnM1Ucsxi73ru+V8psuoAZdpB/YZHQqXJDa54QvK
1mPgKkOFaTvTEn+FY795zaqsaE+1ZjX7cPTuFydaftNepMnp17OflL3teqLavdUfNYK4RKyuRYTU
pHLEsvGDog+F+5RwxesfQbnoS2pTrZelvWsYleUUnLFH8Hrs/M0giotKjBrT98MX7GGS1eaRuq0a
oXjL5ri1nu3uaOK6fIDijq9Nu6pdenn+3HHgt1EqRp1LVo17W7VPHl+7qQVhHMytynoK8MtCN3+R
5oD+dDCrk8WK/MDqW5Rmw8MCs3vXNRlshPt8t/LdCZliS0wB8hZvugmOUmSmPJWUJ2Q7vqLSwTFi
5K7oNO50svRdURzE7Y+BonkdCuoJQaFl6NvnW94tZVV+DIqWiMe+Yq9Pag6wFLqZ3F6RQjOqmeEh
HFtH7Xyy6H4NhuTAL5z3NKjR6UIEXaW8E3dCOkLVhCbIGEBv/ovCXQ4KKQ2WM4P492fFCymksj7t
mAoTo7b9NWkTF2cRio/HmI+CxNVvI8qiRQYVtdTo//uIoJmGgmDqaESQ4n9wcwGiqteObYYRweqS
dSXL+GG2eVp+YQq9ZMV4lbGX14v6XdF/Fjd2g1P9bKueNKsRkkhRkSZ73ZZKjkQW9J0oZUVQd/kM
KclBKQwvS68tEhbFs4/A0cnZ+hVr3QoFp/XNBcGyDhNd3RErfSwWGaW5/L/gv2Fp+ySqwkPpV7om
uvg4u98amgarEP0YztgqdD0PMrQGd6ZV1tNOVJ8Y3eINEY46aVyORute25YHAOIjYM82HL2m4j1m
SAOwc8XCPDxNgKQ5h70qT+x/rCJZBAdaqzpcdL81ete0zK4kwP31yaKajYgMsOQBRK+QNlKkskRI
jBOgItbldCatZH3nDZHu9ajr3n7xrU+zJsw4chfzAkUoYkf9pRTFxFnt3vhyir09qbf7Yw1adOJu
CO40pdM0/mwzd0iG+cOaR7/adoUvfv/MPUIwuJNskdjfb5GZCv3jGRsU8bs9YwXSGlTX9ZX7GjY0
CQ9T02p4DA0EPmb2ZuPScvPaEyDNH5N6LaVD0a1TsIX5YmWz2yIy/0SxaxdwhYV38eAUSRkfzLF/
X1rxxNLH2ZEndZJTSxusVguraQLvZrZGqjiOXbIydrk+rx7RCyA8it0L7Vb1p9NMTR3lixhx5hXp
Zw6bJKlbMoOKdAhmwsosgvlm2Htp8GfE4hTNCVPmItcvT78sLqAcCHEdcXw2i/svBjIOOCJN6TGJ
Di5BWhBStOEZ2VkCZ2MFPI8BSCe4YSetk9XqGrbL3K1ffUnPQmBUad4WNhTy46Jg5s479m1dLrZg
NR1OWWJyfAMVcG1XbFOCabsYJ8jkhZ9askR4w7g+y5oET5Ukp0LE05IEuueyFTjJLqNBSO9BWCsT
KG99NzHTD1ye7R/lr8ghrl+svmfpQ1ZikLuYHrhG2XXJcA5lRdCwFssyB9nf/1t3DxTlIkEq17KH
7XzmDnRr/NL7rkT+YTEYR/8MJltZSs6FP4CJ8gluxzwZuWeNWPGDeGwu7ki6ndILoFe3QAVRN5s9
PdY9rxzh7vmU+NmyEga6Ocq7T0Rg8xgnJJvs2XHrpAUYWv1z0Y7DrlwCL2K+IoGyKHyBtyzN1wuT
76vAObcTZJsaN4MHJX3AFMjG5rq+GF7Mfo7oU6Kq7dpXvLHLQIkw0jVYxpvBAZUe2vBsbKN7iGXB
n65JQhH0FSBJr4VcEcpa6/yz5pUFHogE78UWA+B7G4lybFBYNVWyf4qYoSd2tt2NGw6knEgoDq/L
tecvWJK/skIxdG2erWc6xibrF5LDJTLfyu8QSg/I+Y+Kd09h95dDaMv45gctXyUX2WFdXNHZaVKi
71h8+DiHKL8qTQ6w2MXUbJ7zCikjpDmX4EQufpBe6rshxW9TfNWcRVQo0ohiMRyqvsZ/stQ0+Vn9
sYEyg8+KU4rzj/HBjjsHW9BJrdsydXejq3zgz+05bqWQgOEkfjMwau/4RTGHGeIE7U7IghUSmqml
R2QbyuKPY4jCmYa3t1uCmBZDWWU7ii/boT/PhxeBiNNyjz9qV+jSyyHpjx4CZL2sRFMfaG8t1dDI
zooyAvAd7dgs59foLCe5Y/fSsYO9QXWLuTs80CI5ghC+m8v0c7wAq/Ny96SLt1HRL9YCwId7hhSf
FfO6HlRQrUSxR8xFEKtYws3INEoVpTuaBjLScFTuvnaP46ge5BgCKn4OatB3Orv8PMonO6IeHiXA
0m+sX5/c6zkP9Rdk9Ksg3fZhaMEZHi6OurHOtfSMB/MZSf0n2vqTjO/CzNkUMEpE3wSXzTPp6yl2
WCICFnbf8RGjjaQpYSrFzgwr6K0H0mOw0mqP4mH+EY1p3pmT/HyCX2UtEyaTXLsCMqYD9RqNUSQk
9TnXu6NGWQxGqeaDvNy9eXJtw0Db6GCHFwlzsHrkKDIdSvAa8ATPzYR1pbe+Ywg0REVuQV3nttRB
7NAfK59JfmGP6aT4JsFxgJrhgDeOIazFtoAHhG2J54sM2WouRtVQ4SafIn/p1UU78aBmlX5oKMdY
0cJhqfruZbLezG+edWHYLFVj9K9799N/RTmIQEpR+Yek4yXkwoWavw7IrzcpPkL8LxbsW+rLQizr
7FqaCQMMsZWNG0AeOCaMgEEE+H0LJ8oMXidE+fif+LaPf6fTXsh5GKg4j74tB9OqRnWpV5nfStwC
jC/8Qr3IMlv6WVzGyqomFXChk3DaXZGMB7rBpBkqB4Dr0UH/60V3/IducCslIPJ1+d9eRI073Sr6
0UFKNgAcayhBjPjt0cTC5w5mwzhTOBGtnrepi7p6zC9XScTXMtZ88Rbmcuacj3d+M0rDg22DvmY+
6ymJt93nWeVsFecQWyDpt95ozHbRZNb+FMQqOlODyUZ6FpDG39VkxxmImUdjabBAa2o/eJu2ntYB
tIc2hM78norQG/8zVcu7GbMMCckERxPl2dVrEDI43CcnJrmrRtZleATa7rGu07NE1ApJs5da1SZ0
Jt+cvD48DgxkRotB5re/2ZbOtI+Tq7JghlgHIw2fa1rNA2Fl+eJ0JRoWgfHqNWrXi0avAfoJAiL8
/pGAq7M6GLrro8Wz52SDqI0DmuznrKDwhrOg42BUBlh+5Rj+/P6DZ17GHTjY7SLXU/sb2Qflqhag
F6ZW3BJ98hsN5gLYrwA8pg68Ei8c33m24vfMbnyhCZZivgeLVZ4tPd8Nc4a433/EfeJ9yp4+GosG
c3v0HnoPF4rXk72AtQVhol5zyR8cMdiP54UmmFrq1xYUIlL3v3nSYu8S4nFBarEEnar7ThMZ22VS
GSp/pGXlnAAmMrJIRT9W9VUGq71qC7fq9Ga5BRIGJH1VHxPXuZaUkvHrCQusIwGg+pxdpN48E+V4
S5RG1y+9x9hTjrCFxljiHmUXItpevG2o+Ti7dHwrSvTyaCgyUMNncZWAe3f9UF62Ig5XFBzH2wTV
rfIPyGp7vVjAyRGr8G4LhDHcrDHTur2Gm8m+UQ9Zl2vYODAqaZ7axfBUjXKp84hCfA8nDzha2z8s
7hBylqBZqX2XE+Fy4uhdBag+dJuBW/MzGtc16ecvxHGfasl3Yp4F2xfuHiRETa0zN5NXGeSzdRVN
rnZF9AAju238NsZra2xzWzYoEmsZt8Dltd10/yNIBKL23G/MeTw/ODGdYzIbI4MSUK0EIBMi39XR
Shjf+EDeLVHHzdS3FmifoWt+NlIL4v+E9jk8/PCbnn7HTHHgEAyBq7raYz2Nq2DJgfBMqAQl2JUX
1sJG9V5Gdqq2LP6eKgSVw651Qj6ZG3R+7zqX6Cqh694mxLicMY+sK5aRi2fj9OG62ksqXeHEfzDZ
7dhGTX2y/cCPX1e4BQR3+8HPHI4axGmYTIqJll+allQ1uS+rG7FGsPYFlOme+EyrAc7V6M3mQeqL
J8VbE/9ZoFYY3O3vVkD5To0yS6dny49uJ+JjgwhHFFCq7FQGRklSiIQ00PPgaghyYCXXgZ+l1nT+
sbDIVjW7BIx+lsIgxAbXn+crWlMwCmP++83L/FCbqdIDiQL+8Kvcj2IIEcvndmWWqIZMJR7iCOgS
8Rs3ZbrJEAOJRhMVcUy9F8Xe0nSF4/OFDFQns6PupvHoO5g6DUpF0/OTPoYWHeiRvJ2X6GezY9/f
0mlZ6txqEjenc9B2BHNnVxJiAWSV78E/qUhmIXfXWQAp3sxIiUXk2FtxmRNAvdLwvqtXl1eNmjEI
rVunV73tUi4VzSf4QhazJOOCOenGkbJICGjXqz+g8yJE5+phVtxsIpB8bXYC3potWFBP33Fy7GKr
AktJ++S7tPYmvIvxD25j1Bmm9b7gO5qWhyW1Dy4OJbRPslr75L3wYDKLK461TBgh64dVTYp0DwDz
geFiCh74mYS1EU3QX1kOPVamMi2eAy5TnQ3I2Uey0t6lJMexA4Oa+HYilxKdIekeCny316ZDizfF
KwPtsYs6cm6U3Lm3MqRg5kDpVRuV6OP2MBcosqCwVB1Bx2gO6YU9OJS/YpCAqFDI4st1tQ8Zs3FT
JihQb7ovdGd16Czr0QFr7KwQ2ZtbbzuRscPC7jF51cOU/hLWqC7PurSr+TSkM2OXge2iZTKF40hB
QXyXiSsDL6OqNG5w4gHQpqmZU9wtcAuWtMOG0yUSqCjDSmefXgK4M2WENt8VrJnD+/yf4ad42SXd
i6YYCyEC9gClwXYB8qdoHJZLLvaVJ63ZdsovuntbQSNPmA+aSugTk5fri+tBTGaX0xFrvq37tjJj
m1HpyBGiqf+26gpSYBCA5dOfVrBRVgGGwBm774xhFC6TcA7KmokM3w6jpxzrelLpDB+Sa/e6xnjV
+aIXHtTGzZUPywo9FAV7v5okymddglMSzOe9487zkFUPhcovkmZ56ey35NOgtMIzzby9vSnb5Bhv
n2qvU/Wst+JOzQj0VQ0NTZh+AVIhJBsFRtiwyc433ThhhJXqan7THJM8AsrY0wFYSlPB+P22uaX5
eZusHCwN6X95Sdhemb9D3hspXxzcmxUtwGfSG7oEAxoKKUkQlnkdxwLQn5tEX2Q/EMQrhH/Aya3P
gh44veXhL4pDSxt8J/dMpQZBpASY+WE4QHWJH26zN6diujx4l1ImJgB4BzU2Gs/gTiexrZWKw6WM
Prcs16DsX1iaCwIEJeTUkQBUCCBr4KAk3RyOKujVESteBVpR9LSPT0OI7duh2URFIn/Zy1hfjgQo
sQb8hnXpfkdoJRfYQTGjTHR393aQHu9i3sEU3rfjYkE2fFGzgH8W6uEg8D+lXGowCwy6OPKb+Eqx
wkouvOUNJV0HHjK+rpc2KSmquHvsNX/79WH0Vy+mOJPUH+1BBy03u6E1w5IiSD3UCxx60PnI71IZ
QfaSw0WC8gT2JqYPVgHK17ImJ8DIUcLJfniwXrbiHrl62+ww4tGlNdo2HDS22+s8hau4UkjUsY0D
V+vthoFxvoA3DG/wwNW6+Tx+Iu/d7LvsOxvi2/M7B/nCdTXMQ61279OIlpt5e8Blecjsx8IRiNVM
PcaeTFFvOT0TdTl5pKfampFBVnMePhkrgDDyvTpaRAIB5Fec/nOsHc1JX0Zc+S6vvnL48p3Da0MR
WnDnL5Bh3Fnn4tUhGSpKpUVnbmO3eRPfagHS0nIGibQoUZFmMkYbobzs18brfPaZWutY9R9wso1H
5BcGCHVdjgYB96WZXpLkjQ03Qfta4vQksTnx1po6eMnZvlyESeL0ttQLSwGrS7J7mnjg5KrwMdJw
J7QgzPvBifomSmAe4ahc7cunOpGY3B6whEA56256NALFpQ5vtX0qsM8FEQ5c0JtXjR9W7o44vS1M
KBo3ItJxCODFSzIZSDPmiPWjvs77smdLLZQcxi4OlvyAto7uSQ1GwFuzmY3u/cYN1i8lL2xPaXuo
IVwsNd+CUvI+QC74tOqxwP23Nerw7/Sz93+dxo5feM7CtKRGeIe/WD6A416aXdPWhAFdCWimkJOd
oG7vPsQMn0/D+VkRFZe/ApmgVvNU+Ck6l5/qyTzVH6vPqIlEX2pl/QK55f0k7FzLCkNUJqbjPWnx
2ArqOdHWH9MeP0QRXEnOM7oMzL3lBBpi8U3FSqEbJMHGg/ozD4BX6DRJXXyceQU+UR/JvGVxjfMM
hdFbz+5d8mJFIPFl6QBiFyvAuR6ZbTNnJoxn5Uo8VDFE9MC3bNdRsWyajkpomhEdquTwmdX86GQ9
bF6JStQZOSxqMwQK6xHmGQNG4qmr2s1126jrsfCaptMlZSPcxbuJbaS86isWcnxsuqRqPvgm+kVE
a2w4iYscBmOr5jRFcPfkh6eYORiXqgdUy6ihR+5FM9zGQyCKLEJxqeITapVd1c1iHWx6h5LlbGpk
Ifl/5RZqIFeFWbcJJqzw+3RZfvzI9p8/Bnc2dacIblPRqtzubYfKmKEsoiSVvEA6nEZaPP9dywbd
5v9v3fQR9WhS/rZ6PZKqgIrxFOXyveBkes1nYEzJHbTTOZA0ptcM+mh7Zq5pMRQAJyT/0M5NflE+
h5R8izU7I2ho9k+45zE2iTW7Bwyl1UTKw00GjpODwYmgSNDGCfHNMkGkiFsRwbcXE6OErHB3Yiyx
Gi8wbCoVZsd0cUKvtrS3JVUyTuUwGsynuzE7UJf5oQVjOX/mNJ0Dr3uYpAU9cK9hcCmwzex3jQx3
XRclopUeFQaMJz04fI0Y1icX3V5hwc5kHa9kfD27py/FlQUp8KQUPhnVNygZy1QoOg+EStJ5AQIN
3G7X2uKVTRcJ6yHlUOI6MafirCn3wEahIV3/pYKj+wWImvrQlW4g9DbFrMiGCjc04Jz6HMnnuuZp
WIWGAqgnFv7RdVJnjt5ydpqbmNNZip4ReQLnoB7mAmZGXYAfBv0v68gt6jmjFvmWV6vCXAoo7k+g
DnJ94TW6r1MSIwsMXnGyNE7IhFC8/GxHxP0q43Q0tiosZLfPBtG59pS5DnSO7HRxnXrsB9ir0NJw
7ztbJTpETHKjqgrMqCaK/Co1w9f8O6SisYW1aULCxVRgldFMHp9TQZsA94hbs6u0SBy3F8aP+R5z
527ShtiAptY93qlQFf/e2Xoz8WirNriGC4wCYXIXgKGhXlhvg8+z4jkeJmzuYEN+N+BI0n1Q6VCF
YCwO9fb73kCDu0LMq3LMNMzXWYfiFCqDz1os03jdiSYj5YEI9GZbj1sE1mkRE6NVmVS1Y/QDn3x+
jSorHjaT+c7e1oGXxe2Lpxcb7YuaYZO7nQDTkOd5HY2heDOQsgfGEePLJc+Cto9KE/MoP20MLZSK
bJXxtfNgyEq6E8/KVVLfTBaybjtxJUwDA45sR0qa/SYdl1vaZusNHvAkZHPRaIHceWR0002I6iKM
Nijhsavw9c/p3uNRYXCjaIBy98PuudH6dkuRGAHi4FgvnPbX/46ROrdSYHYqy/b3piZOI8kXx3So
Wj85Ddy2+0vKOElRv8XeOiAGPxs1ulQXthzIB69owawC31UIvHqDB6O4XUbqnaq3OG7UStNE6q4z
ZipYghcUy0FjFgTXt5u0uPBQi3YqnBsBqEkPZF1KBAdkUQPM88gOMe7QjyefLhYv/p1FM4UnZTkM
iaeehd4z6RwdLdFY8K9GZbTcfIj3D/QAulQkUZPDLzVudZbKUPU5LHfxgxKk3sneFesobU5uhB4q
oNsiLiRfgYnSCEYL/JP+JMhJFHg+sqszyML4GOW5hQq1l6qJBMPqrJE89EjMbpKWlWZieYSzgNnK
TMyEahSNkzU0vMC9AAi7/4rjNurYm2QjqJWd/JDFgpuMwzIe+2+JhWA2iAmU3fdSC8OdkpyA9mSJ
nyNTFMG29YEx5DnYC2f4nuWdgg3SKk8M6b/NKkIDVRAM9xx4wPyVgylE0pZFEa2PaqwUhjm5A79L
D/4Xt9kIpxA+XQ+/mY/BhPaa0zuJSEFIfE3YBcEUllsQedKDxV6bKGICP8dCTfEMgzBSQqNXqSls
6CqyWh2MZ4F3wCkM63aAGNmLTy6mqGpzb1WP60lk6tRciH/GN8EeP0YvdCCYPI1r2DI9g9uPVm5r
KThskCO+qeHte/oO9AmsFy6R0YTC11ufIJjTosVyPTTm7B+dYMXwdCDH2ticYbPQ8pC1RAjNj8ct
J+dNFQ5eDGcpurVRWHS5qOuevBFHTXHMr5E90Ga3V8jQSKi8TaBFqEBidCiWFOS6KuQ/KMYLaA3u
aus8dJ3Pc3vbRYzz/N+f2BTt6D2PdZT/hOBuH8zyu3+Xcn0chi+m9/ixP2GGYLVQNR6uZKt6/k1P
EpzLCk8sourbRnbFzU2utoBnAJH6n1UlTE1mcdgxKxnl3mg+z1d2qoxScAVBKJNTQ2q9A+CevwBx
8Z1yuZfezteRUZQk5769qWKvnsYlS6IcwtfI5DQ8i6QuUMjo0V5m93RCTJLJiSlut/9t31Lp9iXY
ZsTIu342JxblMpUnISehpd7SzFibbi0i05NxhFlRYuR9sp/zZFT5cThMcpQE3GihxgGrhU1AMcG/
PL09pUbOE1bzlBHT6MB9fgs8rIRd+U2AyXjDZIibs13CQsxgYvhGsrCRhorv5db/RBfZCfmxXdJt
SECSVG/W609WLOWIAX9CZjYsQ29SXdcj6DXYo+NVByZyXXUocGNQKj4CLgZ0Ek7dmQ84WNpP0sQu
b7m3464B9Wgc5a78Max2n5LvSjrZ+yqR0vQJF6ai1JJe3MP1w93SeE/SO2uK2WVbGP2jKHq1rDVH
Crp2rSYjUa7fU+hx/B7eWYXyacX2H6UgNlBMt73x7FvQyZL23Ce/4Urk6TawbCVyB0RhV2Z1Bghb
LmLM9oNDYkS3h0LtOd8BCFBwcR9WocZWxfew2amSGVHPoFZeeEkpBt4fHW1EL8LZIHyDkKbUpdLt
+0EoU7j3htaeWzJxpUgl94g6bBhEHM4jMjR+FmWglSmKrzo6qu/CpKCEurKrVSYYQ/6XqEF3Vfre
M/avuaoP3wRL5E0/IUS0uOQgs3r6cZmnGstLcH2h6Cv4Y5YnuogkCxxFpRIvjaj5etFVNlnMpZoe
eUzz5Hj+hlGo781jqqRDY7ghHdkN94l19aJVFpZ/EYhT2SAg7o9EdV8/wvx7b8lZ2IfWPSKQmagY
MrmgEx9IPhLkemfl6YI5YDt6eZJeV+zPjy8m1KxddPyR8XbmaHJMmvdMCOH3d6D1ZDxraanA4b++
qJ3jVLry5lFLqkMNt8h43cQd1NKAP/N576yiNau9FVPExnJUQA3FKpWBp32vCiHXt7yazVzYz2rp
0v/z36cpqHespq5zaCxl+v9zedSJ2KTLAIL3aBQZgu2yrM+SURiT330F/mb7pAUUPkw1aejwvmr3
f1wuB41K561Jv+1SqrfLKDvjluyjmjjQcsLUG+VTX+MlvmI7rUoVbigiYA954zZbiS0hokuUUFI1
Lrrwjcmi6uPi1zRH+5bDWazx5gObEdrTd9gwNsgiKYTgn+ZPFxJNjIYs1lvRK1YyxlYJ/WExs/np
oHk+yd6eQKjuqO0KceT2Nbwafz1cDzBFt5cyw8EKAOMyZXqbAuYWZisp1fBGRlfl2FimJFPSwwVX
ejdgzeBzYNOibP2qLafWLaxk5q7OwP8Ksf6BViAECKfe2oYzkG6fh9JwGW+Guv7D5NoFFrEKLKq3
vbiuYjs7leVY0sUpNtbzOGCfbFEuixxoZhyqijCRwQ+tLUjF7wQWNBfS5dN/FtW2IQDSsll1vRdg
nGmS0kg6/O3HQpsj+UytHCBnzqJgWkbFJYxSMH3aHYvAIv8uHQ6Em4zEXbWEgT4SqM5XLIs6lFSQ
V+kveMNMQSUnLnv0U7DH9mZcfAFZ6RFN+9qmszZxXKzwjCRyx8k51LphFO4FcH+IAayJXmLcMEqc
xyfOu3KLhifa67eKM8pc3huVvSs2XJut/IJTx63MAfydWvwtb79Qt5Pq6tWzoyRUeK/evC6jMbwL
Q1T/d8No1cFUKL4NXjRSxQAJO2r8tTAMft0GMqUsD1PT5WuRGJ5ktkRI8RlrOPAyGh0D8/grBndG
/lq1ezc/naPd7mNr503qcw2fMBM1LeiLHDaKEAy+vEdrr7hJdQgnU5FnET+m9Rkj8mxGKQmMOqAH
fDk5Qpux7aVpTXtCKE7zMG5cD3s8y9Dy1tD+7hR154i+crzp5u+emdNDkkf7gJWAv8ynmukRoajE
kg+IyqcKBy0emvGrwfj/g90nqlQ6XXVBeJBx43u2YCOqSo2MiiEo5pseyvptOvU28d3fWhvFfZx6
DWWp5O5dNmyLKy50RWLGzLv7SstiIQhiKoLBJJpwvD9cGkk2ISrLb6QiTtCmJc8YxEqbQjPp4x8p
WNk5sUQ2iCGmyBMxCRR4YjqAo9By9flxWEqdhNBvskeVrKjZ7tFrkPkwO92hcFd6N7/p7/QptYKz
EuWrlDOVBLrgJmKnmh2H3MKWbP9MztWLPoaH921oPjmsAKbSBAtqG6TiagstbRfr81FgUkO8IozT
wUkFPJfrHwOLdM6xsemNd4wc063CBBwLUOW1ucBaHK2CKSLfkmxtEV0Nm3Az6nR4k1UNLvDHaxHs
RiD/bFwNgJeaYFFHThUIy+WSpyti1TNLbavao+fOm6UI6/bXzsj0m6qv3QuC4+hMFaj17bxVUbZS
WHSREqMcKMd7oyjGGaak/iCjvQ4pxRD4RCSObO9aJVZWysfAZ/LPaiGULIwjRz3u2gDccgjzjhBW
9vrf7WYzuKIuGKN1mpijUlR8hz+u85AmtxtTENe64jDmwVMPVBkmUE9BHlcgorGgkTYAuF968a+C
QSsxEICR1IW5vWf13VWmEHNy8iBlCpNuR1DuYDqloSDxhv6BZpOo8CYJkp4oINU96eMUO2Os6miP
OXukLryZ9FYIfMxe076XJcJBMj5SSIVOimPswBQG6N0U290EUaJTTdnJZTO8yjdlab25CwQaSxcg
HySbS7EymWL2I2x0enc7v3HIJOKG7LGCuZVbuKVMdIhZdOr8P9N8gqghfnfiX0MdvzeL3q7jzKAZ
sb5nfnmqvtpGiuZIIXsuEs829aoAitMdKErm0/5JKZ7U8ZI/0QbDuUNnbo2aK8PpGJTDIML1rpUW
4xOHkR67d2y8SYBkhiZXLCIDrTJ9i2sSS/6lxRnWqDBe6f1NnWDmDJlEFysO44WAbdN1RX8DiCvx
fpETFKICNX4gPSjEZ3YuoNjxLCkWzPmlfX6pKiK8eZ0Gs9Rjn8ESPHBnzhNkHQEmIGJ/80XXmOFT
fFWv2/ap4VL3rnSTOv3kADTAfI10Q5ArHrIVY4Y3fTqwxC7jKxzm0F2/SjoJZJTPjyqS2/zvITYo
ErxchlvFtrzguqvdk78cYwf5/sEraYc7WHizSJVK6BkKVjLtsO4yRPsQgNsTOrSoR4SNSz6Hw6rY
oii2tjagf3TMDfC1AIt+9JnfBYpXsuBO3wzVNHOsFgeScaaN8xXOfe81iwsh/XHXoXDl9t07gcln
2lenkprH6lm4Hbty4xKkrOXDviBNp0VXspsqcUUnToYh6SB1LJTSPUku6qpAdhFpf5fZcKjyAHfS
ZShRVwhG6Epd+iQW1Yrsh+FpDrmRBljw0rkzq+Lw81MTFRKiomHuflA40gDeaUn7e6aKBCnb71zI
ufLL9fI+ufy17Ql4IHp1JQ7qLLIZ6mEKYxVf5bWbXbbwVMqYgQSOJN3CspClUqeqmyzIe3FCbH/6
/2ZPKAmZauf9w5+K3eH6SWcT5DWfQUoegF+V1RKq9Wl3dwhjn6RRvU3eNWb2cDWw+nWZfst5xCv/
7eNWcS30sXyppu+7Nkv5pogYDUg/L3M4oAYwCSW4/ZScqQhYmaKLga3jxe/ypTZtUhbHOPdShvbt
edXraCqge+heJMktn4bWPdmBXoGcStEjkm5IzXbSGfXnkFmPsxCZDKU95JEA8Y0paFrsD2oLyuCY
yUs6c0gdHe9WNRhCyAo9VdKwWi7Odkvaq4sXF2LrLxSJ2kzzh9K3Z/PlUVRhEeda+MENIDivfhpR
1RA/qIl3EeULsQ/kmTQz8L2szey8Sz258KFO4wIsmrIqVt2YEkMqiy8lXcfGBjAPqrXY1lFReZW8
H3F/oXwNjjjDBSTAF7qH8jvHlWlEDyAwETgUG8yMEJtzNAWMnEF7YVY6ZaJ/FYd/McHGFEokS3Qa
yYSAWO9ZYmekINfG+PfzZP6ecIK9w2soQcmrY4LkX4FUbriLOFywH2gJnpHtdLBVWO2BaqQR3jEs
Zz3CP8vb1Ek+C4PADTynSHhmPEdEAid45mCpKusoP0uUhWhFeenQV4Hy/IOnrV/8n2IfysXm7Nq+
PwElO2tZrvXTC9yR5dVa56XXUNdB3eKIWx1NvOackeoD8zCGPueyG1nQ4lpz0rrmrkzRWv0IH5VL
r2Oanb/LCKCeHIJ0PJ84YlQyeUbQaMoLqqy/WXo6L4c29pS6HXjUhHsJsFpoXA7DzyCpb5NJEt63
x3D9Y50oUQW0AfzLVj0RjuTlzVBy6wAO2DctJ9OpSNncaqZbZopIqvQvZJR4chKdB/GdHchndzJi
NBQReBmp+GP6VHnnx912KIa9iM3p6bbrwD72y3mdRlui6lUPk1mSYmJc5zY2CXbSjtJ8aM9lQnqT
8IhIIC42W0WrlI8GqzE0JpEPvvetIi4XX2jsOE60ao8UOmP86ziEfuoh0KxkeVpWORTBjC/EsOGV
RFUsC4xNJCIQzlObTg4tzlA5ojXOapGUxtOIRcylR7iMXAKOc0xYwU0MLAr5z4e87978JLx3JH1H
fKHwGct7m+S9GzIxg1HMV3YchUzIHAAP93AbY56nyj1NciXp/iiNrBhpEWAbUKqIdNkUVQqnsVA8
FwbUsxPssCcMPNw6FQf/EOQzP7QZL9XuAwxvGa5gGlEbS1Vk0Yz4PL706/SLO7nGrwj9p5VTaT5S
u2ciJy+Ugpmsx/rqRUeajK5nhF1YTNYX107RxCtNdyC21udVgwC7xFWVcHTnYfcgER6ef08F55g3
nbS+UH/BOGx7YmrwG4FizdAj8IXxqlfg+CwA9JGlC2pdOgoazIo2jALtbq9A3tLhg8ZIB00DOyWC
++G6haDx7MDHPTdiNZClzaddKzwNZD0XooqIeZCwmTwOYI3S0Aj/yJWi4BGeTm8ljVlHU32WNfup
ldw5LDiP2EdwCOQzXE98uq6k8bvwfabC7au4HIYIv8lkCRayIXywr1wMF5H+TJAD7ft0s3vGOvD6
ZR5QVRpiOXyBrv3AFTjH4kg3Hk2Sx5NiYSVxqj9NUG8sG7+OP2C06j6VaqzGrFG+6aWi760obcyR
B7Kdy9J12n+Sl5BzEd3FcHrl0x7s/KXON9E6U27IozE1gLbpcLf5es2pIKcycT7aGg9OHrXJ5Ysp
J4nIqcn/V6v20VMYMgrwj08O9DddMf5nIADdhJ2P6jF2fQ2kOfLETI59BKnF4/EHlNFtwIXtcn15
/ge7p4H0ZWeZrpNsu0fRuwjtYDz0JSpbVxHGjtl4lfJh49zoPlxgjUkbAr+KujmCF5Sv3xsbw+N8
g3v+tx1HLriMYyuhs8S1Ulw8M4L8URGzO+iEgWwNabjriNQGgzMdXEItAepo+BjjuduUO3eKmdOQ
iYCCAkvPXpe5q+Zu4X0YbbhOe7ulMlTb8Y+m5nVcfWNIbPDg2HoTJhAQVK4qnoxIOzVSq2fnZf11
I1HK2z+1n9CJbbvmpvF4zxFXJlTh6zuo3R8drT6CWt7q0WxTWzm1JNVjloxZtsfre2Dg4hGPPOVv
/SADNW1eiAIhJuTjZ+W0Bq21xGMJApcaUw196ciddKhqMLUUXZ8iI0tWw4O1RRrjxDqoTnNpVIPN
nhYx0esQ3lDs0d11ef/fxpLd2lxS1ZLoT4usad91NK+owbZJlNOlRIwYGrvksWwFSPZ/fA0cKWex
lCCoZxqOesg8L494vJDFYb25GEsY3oPo7kzNNNO1sU000l2alUthj4QbwHvLP87OZUz35Sk9GAJ8
xP55joogl8d61zjJg7P8dQzGNmwj9KY440QG69jASG35uQl9IS37wSUFwTwzhb4sZ4WV11Hf5V05
VyoxbiDegGm9Z7AQav7Ov4bAso2rTh7yBNva0pwJT6m/2NrSQ1mZHzjO/GaAQ4UoHw6HhnnA7Z1m
3wHbLSP003hrHuJS3P2dD7d2IlKgFQnlRhFYBP+X5/gTJGguu5nWbzN6NXAPE/R764pqtsXLTLck
y0TFdTse67HkOJiVRt5z67nTkSNYqMqIE3oNrfNCeMNOVfgzK/JV+4SuDCyBhehyxjxtL+6+wvW8
8UIZArwb80lGFf4bayWH0U531l/43hWpnR8qTP8BdynSba+tkYUCW6A6Ycv8MOpvEafWGaTefmVF
ILREb72BQ4C34h+5h20uXoI5vDZVjrUgzCf6uvzAybXC8Aj2SmyqAs7QA0D/kwGE3BlI0wWFi8ul
ru4sFlPBiKD5yG0mOxCT3uVMAff5CCAtGOSU8okv2/3DdpP1Kjbe44JcPqmRkHn5Bxr/bLm8+ach
m9h0OonYTdlWLSTMvfZbRwJq2kMSooPFcpcihxbuUqE5p4RVUFtcYjBTCodJxnGzel99lpikbA2L
8qApo/c3c9yRkjcsNwMswHkyH9qyqLyyLYBLQzS8eddHL7GirZ/jIq3JfCT+AEwtsnmy1qixzMfm
pxlQq7vsQTuXsSatIuUue3O4G7kR/R0BMBC2tN5lktAX7Slb72kETARB9+FkMVG/FwthmDR0+XXu
Mtrs8Lqn2/aoyPei8hv6p1jGEzsaKn1V7R+/9aukHKwRFpHiMEUjvatz1RHF/Rd7jhDuXkeAx3eA
aQWtu5poBVKdB0k5nkyRIUUmeoHi57f7jUxhl5hrhwRYi19jg94R9Nc8yrEt26eNbzZY3wf+Htdx
W/cbcLLdcR6e+BRrHLbJn2g4xMAc3Iv39COhj20BVmc/1Js8exA5O/RWoh4SyzfuGoMlK4RaHGWN
thm1FelFTK60sCZr01QGK0wOAkj6LWwnz/LykjcUT/8fn6YbhvYgcMULlsA9+DRqLXa7TxYLYkJ3
va3pgJ/GdBfpaCABCJqKa6IjFCEVrpDm9WYowofvr1W4POmGJilsqTxwR3Omqkxk+83kYuHbHWCK
t2u0Khttl6UWn67ORz1HlheSRNOu+bEp0DtGKZ+xKeTj+S/3jrZg+i2vb7AGBngW/XyZnaiP7vEV
ga3y0SpwIEF6rR3P9oXqI2SSIE/rZpEDUcVXx16dMJmLmrDOv8NgSwIkT83d2AYhTchj+hqQQ+vA
WB3Ei7IysGKW5sn3yA8UjbLpmJWugulx70y3+Ti/TKbUU/Ncxx//NF1s/6RS28YBs+fLi9YUGpPI
JC/VWDzUBg13J/2tm94fMMldMHjlM09rAW21TYaguIeoXYxhzyx6zkPlYhLKl6ETNTQICuonvug4
+h+h9Royvx+g2MYvmATqWveLoKTDNBNQn1WXx9LAdkXpajT40wxp6VuYr22/vlKig1pK/1naCieQ
o83OUFhsOFjQBVw8/KegmWjnMzsFEwAkMDToVd+02+h4vZRTQd114zyUv4GCPZyRpUUv8P8MJvQu
RdlJZjmuPnMq548vCSVM3jyGnw5VbRP0lgv6SJddLF0+chuB9d2rw8zltRJsEBRaqoQ8hwnffG1t
tGZ+//8L5nQn/J0hBfm8JzJyUsNcJz19b4CYa5/fvrcy5BaaApQQ18YkLpvHjPkx3LE3VAPkMFWZ
5r/KQq9LaKhj/OHTO/BtZKqv/Eir+9He3diZo2nKWEt+1reIZGLvYc4yaZ9FS19Vg0r01FmyVJ4U
sJ7+nekWZH5D9tlLFuNWFUOyUx7LXdep3Ohp/YMzgp0Ug+bGhRxqrHbntgRWiDXoapVKy5X6GITm
witaR9amqrjlSImBwkMrY1GpyWzBAzPqBLeJCMp/ReJmA5Y9rmof4ZB+2rF5u7aNFzG9BJBX77wX
O1eajUPJfwUERZO4G2ryuNz8T6EsYHdNurk98AvEDrvvtnb4o+67/tlopExMOnSa9opIKzb7Tr6x
R4qS5tpZIfpHa94afoRZJdkaHfkakDSBPZV+jDvm4l3k8TtH+emUUKrBlOYSyaXvsG8VltZ1HUhP
pgduyo/2xvCyUXewE0wlhT1ZPkbtkz8zTC6DeX8sr0epnmIp9iKyLQlp6R2sJZ7miq00OfMueKnx
6X3WVa/ZCov194/MHnp4OGWiC6OamtkXnIzi74MQx0VjyxnhKkrrKHFY6w0fsOcGMqams7bBkW//
iw07j7WY6krxC/JuX5h4PX7v0nxrteSsF174uD9wa8+KKv8ZIl9VKof+z0cQaYnAyOKu40C5Z1Sx
Ayn4sQOWq61RPRgiyAMjtAHUcyTpJKmr1aHI5Zh7l2cugALPkfOoI/n7pt3v4WnMof1fTzxZEYJa
6Bq37qNtSeV3PeILzb6InyNKbLOrVKPZFUJtpwsYw2sVDbBGdkFgFQ5w/Hv1yhtK/jrjlpPV55wY
GDWlRWMwDywJu+McLNLb6ADWgHs7bmblGg5ZXWnm6q9fqE2UuF6CLMNabQuDVuMLokRdn2+wCbJc
5AIUdblFgy0ao9xIl0MKo8IXzALJ+FfYUbLte03QfPGzcFnDtwXIcbkX64x1WuqxIbJ3S6vSvDwF
kY7xKeq1rRI218epNdCo/vSq2hzQSVtSLrTTOrRZoLI84DKBu7GXMJgF57Znlwwd1dD1dcYAm2GW
k6lkv9P2Js5LJ0TaLv+u+nDfnXzHQEkKiDAiokOUsmm3YgklhguxmB66y0zcGydamoGLGkAcNAa9
AI/KLJXUK40hCplqz5HLw5xRXyL5KvvsY/BsDWTB8z5ktiwqgyC4rgesyCyghK0TQI2ngC8gi7wG
N+VJ53CDQEHSpXGtc31KzyuuN0aguBjYBrTGeJcT0ggTCVDAkSbpR5cSTOAwWjLbrEQevyEcry5R
ZEJqTk2uoMo7+NvVltyq13pysDemH9pPz57GJGwmGGohDMgLSIkPFCg3tuztBpcenDXUuvraCUhu
ofwCat8ZLsf6eQtkop9jzYx0jGeXewta36y3C+P9uSCNPSJNoGx2/DusLqh0KIR7/HvdNf7STJzC
2AiIAd6IKqkalXn5o79UJNpfqwXpWvB7NHe/3sbvZZw9i2iQH2eOMlEjLEGwGO8HWevM+alWf/oF
Azv/wzyeApn3zauZ37YeCUBm1KUJzWexbcuP6NP1K0TqqrUI1vj8kTBvX9qKrmo9oSS/htskqh+j
DUnLqFmtV7GFfYTT6S4Sbq1E2eUAwvNMhDQeeprOQtSobNyplfqq3LAIOA9bXy1iE74R1JQQfL2F
FqaXdG+1rXLiACfR+sU0tngdROCaBWM0TZu3628tTXhVchT2EGSe0g0BXOWl3KkNOxiDjqY3PzCG
69svkz2dQp6G+S1yLdwSK8fSM4fWxU6cvifyPq3teI6JXKeCniGepKm+z/3qI7/lXF3w+smD1E7M
0mVuMJs4+ZOImMEKHan4moQoKXkbaa2X/ay7VrngzlHfb8wXYnY2mWBhoPW0NcdiCSHU7McHbZjt
V5Ss5MCuimjnvj3lzD+HkH9hsycTUP30LU6uOT4QfnFGTMuSbfGOp38UcXDpvRiDg2hAhoJUk78+
t03v04g0k30g9PmicEFL9ckJe+13eO4mE0OWneJAudvCwLK7jWHrjYtaqT710M4yjET2yklrqsEf
g8d9qcnPxZbM/PhscP9rp/mjIvg+c49o8qpGhNSsPhiZFTtBdrTY6qnKlpB0rch+mZujnrURJd7w
b/j3cO4Ct3fHLYhUDRy2RRCYakFwOJZ0jC8zZYSaVUPAXU4klIiOyXv++M4AD5Jn8Q8qGdKZozv2
tjQuAWcTbGG7QQlfcBOUtYBpbiz8AjgPtpAiCGFDQwFod64TyI+PTjHGxoDl+Q/6qmKnngRsMtZR
hug+Jc93Z+vyccEBhD1BlLm/q2Mmqr0iOo9APVqsnRtvcZAmVCPUteMCes8d92xKHXTCPanqLxtq
PT85LQ2eTJg8F9FH/ri47WmvSogfM10tZqIZfIQZsNyl13/9++3DRrGqPGhb316p6T1ZNkmEUjNs
HqiIRSIwhzFnXiOk0JLHOAlcbb5EvM1LLHtWOQqUJTBSb8andJqvi6FaH2pseXXgLVIdpVAynChJ
yOl/+83F8gdI6AwSG821bsh/uKap3wONy+xO2b+vJObpvdTnDxBUEg/fRSWqG06OcL/Y6hG12imr
xVenJ1Drk6EMsICkgL4g8vlEbhFFpG+JgCdnED9Pr1EuZZe/q14wYqY29lVDWzsMF093iSWel1vL
rdaqLyoHF/EzecNOpcjgkplkT2idD9jvZgjUL5mmCzGW+Zi6USkX5CcNGrlfaN3gz6lZoEFT5eDZ
20wvFb2S4Wrn+pvRH0j7kaUaBUmBHMmCdqyq4KAvcZMxQ0MEsVvx7BXEeRwISHnx4ft0ualGtclZ
nMrKq2E4hM3N7vMBmq0ITqP35J+4aFxDIVMEvKx9VuBgrLY0Gc/S4ERkPqDv8t7jSi40Ox8sCL8z
8e0n4x0XbCUPl+b3FvcNB/sMm3LZXiQqlVIGQQvoSLKxknmoQwU7xmy66v7h4afiMzmQtrl6Zayv
Nqp2de1doJZhgNQNVF87kcMPWpZqG75Cfty9CntTsxDHL2VVJPB5Z6T5dZIJ+7jmDq9WGWXCuhsy
JVDkCq2feDWCgpEVkY32SBnGZoEJRn6Bv6K7WOb4WQOM+ioHWBflIlS60cu2WVc+aRz9EFbnSQqd
FwW/XSHSY8o+Z+utuZLdy+hcD+jFOGSDaluLcOI1jAzfXdwO5CwN7vRizYlBMQXxinCDf3zEoNgd
7UKltDmZSI7HQUhH8r0+XRBGkiJjqJ3EiYZRTV7plc9hRmW1G97xOG3hJv9eSYS3rvPR2SzT2kVT
TPMEJrq5Mw1KLU/GXzVxdY3vKReYxivZLgafm9AtM5M/k52Kw5ZH6xtNdumfpGJJx09jDVVDKC+w
4Jfn0Xs/g9r0rOJEhSmqgqXUxQVIcDKqhgFpdGai2jLhgPHZUTpoQh1s67K38V9kg0gdDhVM6Bvc
HRx9bXMY2dEMcHxr5RtDaBSoBvmMRIcqCKjAPHKStSHtvBTdrvxWHqP6loSJJNfE/7OCRC+blD/z
7T84YG5jLcPbPWyS/h52+Th6YBIZXa9u8cmxhnXR1JCJmBuOalFEWHsetopMSPmYQpc6v72nzfxU
aBaBlVKulhhgSQt0169yHlDeVNc/lY2hVcCeB/mV1DWWoIbwWXURO5U1cEEoRUSJhFtjWy935Mv8
K+58T39LmvQKo2ZMv2zJpfJb2rY1+T7lgYfD2yUPBchBz2+ho98W2p+1ckwM0mcrh12QYgH79buN
pZ0WfQlwHLEyt/ylQwX4OXMwTAxkTEpQ6sslqSmIRhVJmexlkGivLU35xcBFC5Z76vuJeqIKcpEW
o/IEVL2OsDMuQsKybQHmeR8dBnzQbwL2rzzVu2QeaiyDFl6b36LtCKjv6p0oJFwKR0j4YbnyAmca
CqkQIb0oO2eEHsvAtuc2Bin76YSIW9NjFaZmA/LlTJBA/p3pdzBO3sMVSuLNOXmjB6BEG3cFLoCS
muaRNGBvx2ubIQz5+wALs8pvjn3CGSkSKvxyhcXjjFxEGrVsBng3t/SRi9JCTvf0aYsQx01WQWYM
NfRGVHWySiC4IRBneO7hhVUwww/5Hl1S0AZOT2uATwLsaxvV6Cdy9Fr/wZWujQjmAtnJITvPNW9M
WtT0g4cOmQpOxXuF4oX5RnY7w/vH2BYkQn8cBzLMlE2XxZPKYLs6yGS91cG3lYNSWzsdaU5WM+5b
zKap99Lbplwft01wYzDChohbDUnTvTgI+cCgQosogyvnUoUFenoCpr+oDJ7scyVQ/2vibl/zHhYW
8b6supsF4cOI5KLgjsde0MgGB55Fava7vnSgmmtomwtsYDcR2+OyLffVY4JXOX1Kq+uvb48wbQqy
5+d4Ml4zjcU38UUr6kQlNV5Hp8XfBehms60tCHHBhEuFLxF1jXyJacTQz/dhUCFH1d8NxCoYn2Z1
46sBog0M9BdpJ5mRL32J5gLevZSnXSQQDtKEkd/UFwB4TrmXSajyVCGeRTXf1f83SdfDa6M0W/4H
wwLXHAh4qG6rIx+2R2Etz0YbB4KHCEOzdoH/TW+5X3EtIpyjkVYxtTQ7rMOE4YyzCdoT2T0+CUoQ
Rv2qMnPfu8GP/+3GZNeBNgKctKlxBwap/pGxyjf6jZzNYLTiQvrE5JDE8mczjcEUyZCxgqaN3ajN
taiMcwNwaXtQG61eGiy6VvoW4Ook0xPGMJ0B3LFGC2H+cpUAzfeKeR7XUTMrok4vgOw49H9teeWZ
sGzLthZUomzDtrjjdswy654iCfsUVqJ/hkz3VeDBJjcmqC6sU92tfK/QIPgB1cg1VvIgtmVwhzsh
jWxHpcLMzZpll3eqmUFl0zNvOq1fDh45s8Zw3e66T/wDHaGWAco0crHOR39G6Fnpv56boQq1pnhs
90Vfq3ZHihFAt1AQDcZBdrbqDckG7Py784DqDrJ0RBRi3RFC1DY9/5EyT6TlRWImkjlqkv2H0dhg
RW9qdQV2kwU5vH6mYpMFmdi3HR4g/Qe46LJ1ys4OsRCkmUTDY8aHjkpwWRh36dEAv2eU6oGkLk/h
AZdAqV3RPzHWoD7kwXf5p2j0pkmIvt5kZ7ZbmKt0RSgcjU6IqcZI024tHeShD5ZV/t1qmmdv6Otm
VX4LPxaSeg4zSs8fNMQdKN6q92c3w1pN8iAq5+++YBddL5Fj8rPSGaaqjBz8Kw4l85xZ7amak3se
CJLMTTjJGBCfejXolGqQJ7Di2t7oKEDqGPb4I+W1OufLqkOsKGI7hQUcSytOMDAfJjkfUsgudQ9s
nrnFT40jo1J/LLiYWmcngZ88TRumJxUVZv785P0STodFyye056o3oofVWLeiiwJXW3paqlP6iQ8e
H1QC5kfk5qN7CxturoLx9tKwgBm0aci4abe9HziJg7hNMZ2W7ASyHHs6OlHCLG7XDfmvCDQHY3at
HOzM8yWnSE/YVFID68VMFS3sM/DsXXxQJ+kWHtjhBssyyY7h4LErGdBzMWjWXhj9Jh3kNzgc7426
wBfuMNndfcQLtczDgdNuYw4L+KEBC9OPkmFerDkXHIAQiijsb+HOfd/JsuKfKb+gOT+BiEwORXu1
710i6iDcz+guZj/q48bF4nW+hnV3gvMPn0i9Tu9qtxUeg8LNjY4J54x35GirE6BcWQ0sXP+dhcUo
9pVAURqAUD5raTmYs8yMIU37+Sg6E0koE5emJ6GydCD1wfoPMOn0Lm/Hb3bZPnYVctrQ/z/+rFQZ
z2WDDOqDcfmy1dwyaVftpoFJDQ9rpRZSjKcbNJYHWTGFLNzf8txbQu3zArWbgXhAYSRN9ezytZ2a
dkS1/g6rh3iLMr/nFzQVAMupkTHgzinmUBkGscKLZIx1G112v/Qs6mPfiA6gUeMLfljr/WP9mPK2
1f4vxLitvg2i/SXYdSFVXRWoBbpsjmsYMFJEgiLTO9xqza1pbSqTQU+tjeDcxQcg/hRKCMjoOdbb
5Alt76C4C2LznZgknPFb1pGTpw2IuN22/sUxaCZPsewhbsoP5cpMboQt3WihW25e6fLYrbeCexR1
SgYUactkNUkkkVzPR0KyX+WZfllatOJD1MmTkcpz1zJShnKCMLGVBDWsklhvXIfUUd6yMali85Hr
oU7hlc7dwpDWf4gJgH4uGJ97g1Wi8zZFRCslMwu+kHwGcUPBOtDyZQhcJgT6rIeN4UErpYj9Y4eB
vKXlXK+A582vuQYN5Pk5xJMAqjw/M1UONkXOjlmpUIMmEJ1p+oxAENO4XgCIFruzBSS2ztf2a/jM
hrepdkPg6RBgYZ+A/czmUZzmF+2gUWtofpdkAaK3yk7TGrYSv7AyNcc7JcfJ6gh6qSyip0XgMSCt
UhDYKj4D8Dl3eyo6x8r90u26EZABT2EJGSEzWxlTsBAeV3mWCZv4uU+BRcMHOh5V7TmDwawaq78n
upxQPsanPfQL4NCLpcnZqbOed/lZd8o4WIpTSIcL17ookeASNCJuzIQLY75JeXCsatW7BGFNr24g
pHT9AnPNny33YPOFLNMDpxead9obFhVZCE2oC8e+PQuZI/XWA/AhDXzut3m5j1BSrAwGBNbnlDCt
Z15chdNNX4vR79AmsbrfwroPAb6n7oaJoV1Zqxu8+LJz4JXBUcE4tZLRXfedjcgPL5ImaQ3TTZqD
3QS6oRYovF5dJ6a32mt/GuOc544u87Fk5K8lw/bpNac4Gi/popF68YEMGBOLf/OQoE4TOg1pnZYA
sqPG6HbkXn1x2qVoe4fAz/Wl4duTSOY/ntQ6FSQ8ciDmYbD8kt8Uz5KwPbgb/jiYhGNtuJ8kJeAH
FwQafX0+MxFOiMysV96wy0sJ+nftNRzCCyzsJhJqt/fSyCkoQCM1lm/XmD3aJuzuN94C2sQMIyDx
RPjw7nrN+oAckCVAO865hzg1oGCpC4KcXanoc+zCHsqQKqvfqWgg76484mGKKusF46tBHovOrIw3
CWYw8Hl1suHZlFS6eiM9j16NFDg+rhzzdzrAfLNyRPY1vxfXTGRqkJZmCmeWnQYm1/668O3vkgBq
joOkLeqdGGIFGsIy2xxdBVZm7lTh7ddxU//XuxGZf+S13c7WgzEpQQMc/xBShRmDJWxWBShJYrFW
ybQHVH8D5Y2flBxTKRGy11zHGltfkGCTELP5cNGx5FAKwJ0yupxyRYBxKflrB6WXsrJ47qDeGmSD
X0wo8A7BVJ0Hkbf0HKad+mkGxXorUqJC5smiaTTufFd4+caS8KJCkqunoE3t8KitG+EhKOXtWEnF
oc7mz61cZj8RYNndEiSO2CZI/M8StJGs3lcBbFu4w6C37bTfFr2tk4WmEV2yjt7KulMmdM1rGTR7
tMjGPagZ7JShKMix7muoGYibNai6teEXQxOQ/3X8VgqY0KhtCLqAev/0/L+F/J+iIWBEOkxRNzHm
cNmkyiV9O39Uz8C5wsQv3UntNn33SnbGBBSu+UyGt2gg+iF81jkfgc3g90PCPH4H2um4ulcnBYv1
l4gXdkn1Zqaq85ihF0OSB1FindxzHdB5CopavNXue5Nr9PEqFnlu+qoQlWvFlzXh24O2QsOMK40r
FTHtpU3eiu5L6cFnFfi+Px5gFaBFtPQJ9MJ/xKQLj0xBlDnL8chRD938EA3EijK2ZL+z6tvz2ep8
EpXk574yHPkOpY6ze8fM3IoKH25mZbZGL/0SmER2u9nAOlCYnvrdYlz9aEtt2ppS1jDQVCNigCsv
l0bJORjkdMnKdhDUWYRHO5Wp6aQ0ZnQySUJCXEA5GI4ycfrqwIsr1GPi4PgQq2osG/FFVhGiYHLJ
aezZkKhVJYSWSfMKe+8uh7Pt7TGD40ky3YeI2YTxDOemo6yGURKZr+MZMyFkx9TGAGx0P45IvYAb
JhJmWu59ULTbIWBEWt/fMxzE6rKxTbcLfe0ezw+HfRec7nWM0OQAWByV3VmQTHKOiBz+csZyURfo
IGyf+FeOBHAL5pNioOWNjQzJVNhU7FLswbSFCgONDNR+iiLB+rYwzlXXonDp0oJf8byyX0OF/5Xz
Zl5pkOYFevKOzlWJOtGEmgj2pfKorTad7zlrLCFJ+pQ2cV9tCAHL3pJktpRtZavcw3Vhk0PTHUQ4
Eoz2qzSq4Z/Mykk0vie9mlVVoaCo9KE6BdNwewg+NfYcGOkNVxnft0CYUP45JnFrNKpP9MUgqv2a
MXiaUUyGKeSa42UQs/Piz9XdvgbpVBdICH9PB0yjFGYTgQk2xDs0Af6zsn9FiE4a9aVkcZPVvkuY
In+sHIYqh3BkXYc9zHaCFO1yysOZza3b/9TEEggQR66omKukq0AUPqWn7Z5w8B6JhX/waEXFdyjc
69nGnuV2L8sxHgcmbt+SS1U50K9IsaD2u/tNznhY95YSODm14A+WDhQn04+vYBWQdXZvRqS/C824
rV5VykJzEUavf5lseRhbZErhjiZfGL0l3wMh/Qp/bj1mJNBwTuJ7dbXKCwyre0kFdJgFVcyqLV1M
+k4FW209UDzrojowSCQ0jcQrHwRE61QYnNE8MwtyRhTYumugALYh/AIrIW+2KL+CGIVP6ObuP7Kw
lJ8wuNjDEimXu/a4G+LQWktwXHcYLN3Lmpj3BRLguL/MaSNm1TCRo7GtPTtsUy8Aa9aEeUbmRaMC
bvTAVRxCn/k+sZ0Qr/DVfAE3u92tnG7TIOtd25b8T/atdYh9quB1ib+gYVFaj/S+ewuB6y+I6RBN
/NKAy8QBfiBID7vkO35vdM33QsIj2pNVd6olsPHIktZTBBXA+iwf3a4Oiv3uHgWYekuFFy4lw7u5
NjCs8eydgBi3SiQ2/My2az0f1JIafyKNrecBUysBolb7V+gOZWOlKp91d+nPtHAtAMZaILpk+wMU
jBJEucG0dM+gP43Mb5Nbm9/+i7sXuToEq/AZmheLLiLyPJXpXRYVmgdjJDFIzypAMIc1nHio1gGD
sw7XkFKQ4h9+uSm3C+0vXycxgCfTOpDktNlqBccJgDmy0xsOLM57jRhtnNnvJ/hAVbioXYP9Vqej
ZLCGNO9XUi4M9p7ypGzOHdxt03CNNAogN5PewhvJBK7f1hcQgU3jqjg/Pv0bRqdJoxRHsdOKWdpR
y/7S63++bj6KRedFhz4VzKqen8I5eLWIrOwmVqyc0riXmrI0k7OpRbDRGUr0OGwCtVS59Me0iaQu
urxqO/oj2vCvS4ZzyHCzrpnbbWWs47fuFGQhOdP+f49QapZDCbMXVuQrcsHiSpS29giA5WSjl9qm
pzruzEvLBWMVnnHPDTbp/e3r7771x1QJjTNyUI8577ocU0y1TNgQnYd6FU0XohR7eDxY10HhfjVU
qEXACEGQfwYcuZoblRRtv7DL4vtQA+ZJuQXdyfFDWM7bY8k/7t00CDiRoDpVTpOKjcQbLtHGaIvd
6ETkCluGx0Mg3exOsloKoBZvxWrhKDDRBIPiwsKxagAxl5Wpyq4UGn9t2SsldaFgST2qqa89rSeS
pfhlSq0WbBD/852ruQF5/VMeywdjQ4OixH25l+JD9stGkq5u+Wufa6B9gi32DgK18i/HR785kTY0
ur82PS6aBkxED+DZpwd1a/GxKQzFU/I8xdN0VTjrnajnR0DYdoYHPhpEuEkiDGkdgIV1+yh2C8YB
leHu4vZLUyULxZxrVcOj7ZtVE3mPnor+QaMbVfW1NX6GRbMWY8bOQE6QlJIk0T2mbuGbWOWJkKIn
2JNElAQcCQ/c0uEyzhL8ndkEgqrGu1IkNr4FyycByCS3xZUWzkFzS7NJNkk6dVnfI0uzj8n8F+7F
sGnMLgfcnpiXk/UhGM5dTyP3BRKGObd+xLmge5KqnO2bNj2nhfPU1Ev31rlfXd42wxicUfV2AH4h
406/bHDJsjYqGb2CXjcViQHxa1CpP3VOFHAGHMyRUJ91fF7OqHgjgB48eaP/FGQoKWYuWK+r6q5Y
oNQfVb7OEiKyMoAR91XYwSKFwxacy1ArIOhxwXRckqoSqYPB8PR72x6eE3jmxsw6D+RcrHUvejhD
OCse67B1rqRLW8yOieJX6XpQL2C/KuohidgfJVBurJ6BoHW9M3XqX2sT49KVKYrahZx/QMDWmdy1
ga/7ZQu0n8mMo/lJuKRvpvSH1rtRPYyOxqWBBNPRvEZUCBLawEirGvBeXwZPMd7ezn8WgqDBkSU6
EuR56SXiafs/pFx6ConHl1Dm/9UqhXyrW80Jx1lS88IVMBHWKD2fsCtxBdoOsUhTs5OzX/PkMhY6
3Gh/uMt6MOz58UuNfvX3wnZ8omv8Mnkb774HY6cUMt77vQ5HbVTKVPC7Bj3JNDmI0yRh5woScMRF
JUHOUePpuuzDmsy51fB5QkvvMeA4FO0Aso+UOEhBgWASmietqgORDfk6Y2/oC/f9kHGwhBzXug5m
cDIyF+vn0fIj7+8V22+o0sjU2vsfFSAsl30eOuERdXVM02l+jkTry3g/zBB2ODWO1AJbwpzF/4Yh
yn/LlEuDTbuqU4MQLvgcGCV7GESRzOJOGT8pPtJBvxd8DrP9YTpGziV7+9+632uyJfIdNkJVTxIh
yCR1P8/cTipL7M62wTM/yrSdBhHVQFJOba+rI40HMO02XMNtl76sfYBqdTIhYNCS+nvUJW2DmEV8
V7quhW4ZTBs/jPpsx87qKXg4p/lG6vxc835qYqxVttji0c/KmLwSyScmn+2gTCPU7BjgMRNC06nZ
yJ5ISJo7IfhmE/9+zWLmAnT1jwE8VGNvmn2PbcqIR6aX4k0a5nuJmM5ZDMapqlN4/lN/wsDrmi1y
DL30URIMcqGpw8zN8juwT9vpIS86/ph4dwfufQoeH2UYFmUxL7DR/vFUXfSJR6ADU1et4+owx3ly
miEItqAyzMJI8d9nULQXNe9bzhQ7Z8B2hA5NUiJfh+siC2ZoONSuOKkNyVg1qsxzXDEQeEpqQqiO
hm3ASFUcBkwX3528o3yKFSAoyvH4L/ZCklSKj6ZxMGeTg6as0Gn5fTABOQQ5DuAc30lc28Mz2II3
g2SaCJ1ZAbaKf2cp32zwdcaLsmEPNKhHVfPPUk8Dk9SY/ov6eHxLDr3cLLJkbM7LnhgJkasIt7wI
vyt/ppYL4Igy+T6Fu4BlVnzro6q4q2BkI1Zd3u80yqjfPepBzVyesyQT2aAAHbFukism9P6rngZN
LV7SJfaQxeEKLvVp0AXvV56C8TqZ3L/W/IXdS59udQZxWS/Lul0R5hHszeT1LLO6GxMtXslKBlyQ
klW6e+fnhzS8is77qSW+RV1PCKzRg1Cj0swgZeoAzr2tAWV3NC8DX5kNYSyuypkNmfJUgMk1sf9C
NZsx20GXEP+buARaEEh6PrMBKVk5E1ROR4v2DPkeZrSVQCknr6PUZahsOuVhEDWgAVLN6eF3raXn
r8djNpBY4PSaKKgfoVMvpFgbFSMZLmMwPOflP92iSqT9yB7JRvPp/rnFVvnsxaNeNkJl0QH4BhI7
NzxFT8iR2QR4FJ7WDNixaSAjsFrW3FyVsWuaelkTEZXxfGN3fXErkVzZObukO6+ABICsMDwtU0qU
KZkJeaKzOhMl8VsBtxYtuQYS4cVePN47oSFV5qAVfzNSox3johmsSUSkd2vQbV+by0+HGO0IHS63
dYyb8xubvX/BIJFisqQb1PCpDYQtyIGH+IB7h5lPlrKT1U8y5iQxgTH2NtkQwGZ9Yo6GxX6LXnrU
H9xktZlim3UEhrK7h3Lyasv69JIiz7EqJICDcqvYfMgVJ+ElH1qQbLLZyxEr0yxN7OGFp649VOYF
F+8GJIdMYoWHRo4NhUfe06M/8wx+/1nPBKDjZgGRq2l5GIOg4vrHxjjoA0X0DFBeqMiHIrc/ivS0
mdW+b2WrgVs27r7reV4BCAUMS7Vcqa0IW+MbIOY4SCxqIOTmhtvr+WfSBS4Wbr1FFewrW+LeRgsv
QXLH+9aLufI51GCTUCvBLut+i8Yt1eqhRIzRg35vvbG1GIM4yQ+LKfc9S1vJoPFRpef1UCR221JN
67wQpCIh/hQTgmprruJrecEAaWKKdKQ+cwI9AKCZMacMvqxuWBf4HBwyRG/Dovbk2y8dpc1YYbSJ
0h26NNFxX8FXSqgyX7VjNLbbtidr7eiBIsVRAZzd4oV5TQMWvXPfcBPty0VsAC4RvaX0QSVAzN7I
zzC179P/NLlNzCCr5RDgkTWpzGbuSL7ZwCPqBcBHaPyKqZHKjVESQ1Ugyiy4wp3I+wxWyrJBLnjG
2BNJADRXc2g7wNpEiotR/+xNmPH/UQa3bVVlCs5CRSE7gtmI/XGnhDn48Jm2jjAHY84hVZMOBL3D
PGPXSfEoLQAtMfJnumr0hye1izV2I/NvrqUed1sZOeLqn0qo8gG8BZDiol0o5/46HafpopT8aeuZ
XJ8XIIeu7ggKsmZgRYVmAG8mU8/T8GASrlutw7XVCkRGPPr5dyjGwDl66Elf+4AJpJvctSylNfwH
tEd6dBvr5gpaQ4fkTPG3FYF7qjzc1nnFK2K0GGwFP+DAVcsCRr4UT6jDbiC5W0fV6s1PJARy6T2v
4vUgIuFZEd3RtFAyBzvr+dHnhVTex40WrU0zwC1CrzsIWFVW3yMzi+Xsp4hUxTmL4YCn/hc/7zJw
S6rPlHwMVZ2zY6wNf46wkL96Q1i5FwSmRNyYOQfVV8QjSTrCSCtSm0woL8+W+qjscNd96ROEL/o0
UfEs21PoHcaEkHDDjfzrF6oa1HN7wk5i3nB8g+gtQ1s8FT4ZVHEM0QGCH93t98EsJPrIUyevK79T
JjO1ZlgPNqk3psRA62Z8ZInJEVOCpq/BOu4HGzTy/Qiaj8FeRnlR5qpr2Z2kZ7Tj7eFBQ8HcpOj3
mtO0jD4oOKevJPheNadjLn+GfNFe2eCUHlBlwcfcc7yx3VbQl8s5wdGR9p2hSD8F511MSjQTJCqN
BOH95qXhhZyOkhpE+RH8Z8Ks803gxTIud3eSkrXjS4DwGv0qCVvAWEg6jZYQPQM5fDCzrWrao+sW
XrV+Vwa+nG8iDX6K5LoZjctifIPchCGLAFnEocPZgY6rzhF7j7A/qSQTFwUGez+e47vmdooCaPGp
et0qXFc8eb1AjzF9m7GCFXd0HFr/Iw4hrF3FjoBQb4+C8cFzPnAfQ1/GcmDZ0PRndbmC96nxdMa4
nsnLkSODhVFoeC/bTy8Ahn33IaIRZFxNTuT/ODSzGLdcmPsntO3s/xrdOVdXbWAeNK+oDU6DpdkY
gBPxaVPQxq4+cvvRVjhi6zMe+JOgII9HRr1WakaRLCGCNkZLl0sRKupqtDOSpd/Zgn4eun1T0Dgl
6LN97O0h1xop0A92aT5piVdx2fozUqdH6ph7/5Jn3d+qOi8RJcA8ypw0qPrYPJil1zffvpVUmdrz
L0JwAr5o9mA/Wd1VXHiKc/CsYexlqjtNhPWo1cH7rDaaJayg9lTah7de8jCe7yQs1RwX9h3ZqbBS
cahfrXiJ1xNBOI33cY75SgOt2aqvrvA3X91Ta0iDvPQeC0U/QAqjd0RCIQEyqB5EQlPjn8MxTPMU
sZo8Z+vIeg05l5OJ5nm34Y2zcqStxHqsEB0sdq5t+KgiVAas7T8abeAa8PsRkR0I6LiyBGaoDJcb
2mpskNdZJ5qFk+DENv8qCf1SkXCGBOeohisxd/33Tv54Wsr8nNIBG24ydQlvIiLH0AnYoOlAFu3x
Yo+lclslg9gZ3Q3U/3qjahKDkZ7aL7hq3q85BbcuCcibQJq+lRlmcrwizGGdcn7pzzWe67T1VHD7
UPHjBr8SJThBgUcVGAViYUuegbU56CtyTdrEnke45QBPlu385bekDfNmE5Io5wnuKTfCwWNDPfeo
dNSh8UdOH5ltHf49PbTb8f0CeYgQtqhBr7rsRda5mCptTRUhCsTTq4LZ55aUvuPgb42rcIyMiOtk
XAGGgDm8zN0gKQiqOuqlwK31v1UaWnzbElmYNaofKdb44fbDmvyONbYpBFGsU51ZIkEWoqeJgFi6
2VwKh+zuWsWv6ZxzIOYMoeRdL1cpYnaCdYLUyGUTp8dSzF0TPNPPBz+dtjVtYkWUrCTBOgF5RC4F
UchMK/pxFo4RvlDxbUClkvu7vuTPoBNVyyrko9dmBmCOJ53LrJuPate+COvMzoH1eI9nQZmwKWJK
8821EknKH6xuDKtJQYKcwGlDQfmR0ybVDET2CV/w1dHpdswrZ96q4Aan+c8cUjeDZIje2zSKa/K8
RlQVc50G7stSxaoUUhlHMVoWG8SoAuSfEhv4gbYQ2g18AmRO0obyP6JOwniiikUrgukvicY8d0A3
XaJCXIvAYWSN8ObR/7YwfgtUxTcxPoBbIJqlmnSLuWTxWlJdaftuViH2/eyXdwYpiZyYlu1WyKZS
zWLufMLDSC34OUDx2pEyQ7wqFObc5hgbKrBZwr8oep8DnWBF/KDPHCO8UW636ssvmBm+RVvpqEGP
JD7+B4WVptMS4eymD+Wk0ehzk+xOuM1tUEgpuzxWxzONBY2X7C6zL5Gc5LebQw1YlA9DEyY9Rqgw
cB0rm/gVgpiGqu42iGJsSwxRoHlkfsuCY5XFPmbEqk982yw8/1k/cBzQGtMr1505LyXzC892CqXj
pzsIXrkJCqbic5Xhr5F+IejZSRxt3mAQpe6mFNL5tMWDE8VqVmjnsj0TlQSXEVFiLm0Ga2N7+HkS
nZYRUZiuYq/XKUzySASmeNO3gSEO5ekuV4ib9pxBt0OMs/NcHQG2H57oqGPrIGmkwQ+cA4Sqke3m
/dvwlt1PflklCJjjQ+L3gAM3TOlKPgAMJFElOTwAqLRSbRg++DwWUGKLAbchEGXaBACSoG39nwBK
i+t3NGj1rJu/NT2MJKoAG5o38VNapXcnDfdRwjJvTwl6vhhgjMO932c3oHVHLXPZQbLFDhu+WXpd
gqeoqbJ5/WOJBkrPt0gr+dqgbMgp/58IO3/+CyRs7Hs9iElBGKnEntDtssauDj1LtlQsZ+/f6nBL
XqWi0NUl4jJmtgor+ZL+CLtO0rSuOmblUCQNy18h2Zjy64zBMUkT7gxgzUlXzIZG1RF2gTN/Xl2d
22fMhm0hxbAS0ceq8l1EGPe9w45mJGDXtMNIIO4FSz2s61UktWFWFMw1FPjvhPsJazxqMjReWK68
DYfFML/C187DAfln2i7Cxaj4a9Hicr4GTIYxCNh9FwRa18T857W0w94MHneA2yo8JnsQrcYpt7Vj
UaqLVlx5j8REzx8mZabnjPtIxZ/uydr7O4tXVHmkit4D5mlGKb1kOtrvJkNJdGzNOEDSjjKyHGy9
YvgdX+C+AHHxmemxjxAavDEk+f9LksID44f/SLWn2JZLBVZC+GxHgQD9yNZpUxEqH1lffuKzvmWt
KcpTbLxQ1VoqJHgq4WIwYHtqcK+6wKWM2Bj74tzs7JKeVRYDlbt4ZnqPd72pvtFwHOaITmzJP/1P
KPxWtUHZ4e0TRjYPTAd93wSX/WQqEomV5aQObOPRVztOSItslkBQxIU2xC5YKS51iccktaNhQqJP
DTcEM5aVd/xmSLpK74aRwZV74mqjNeKRp7yBWdMeykV0MHtsjQrszkXpAbr8K96MIXWjIOm2YqwW
oJ+F4OEm0RgY7hQtKWH8Lf2Ey3EXiJo6m9aJH4D/3/gVVFToNNkQzutkQZsByz0V5JJ3YyTULXKK
AnET6jyHNhSJqnISHpI8OckWNU1H2pSb3zx/fpI9N/Evb3ldnJ2IV7Wpw7Bg/4S7vNWzujDUItTN
oRyEhtARCkbuOo37Gw83GlglbqrlKQ6pAogTjKXvrGXy3y9Rbc1aKt+uEJhpQRpuVYDtPqfasy21
ZKYEZs6AdAV32jgPcVwpDcX8YITVE8HF/UssVN2beL/TK0ykA2uTieUhKF2nhmN3/hrWGjbyRsXG
PTzUQGBPylk5jCc8yU5/BpZZ6cGqoR2Ya0o0zHXSVzCVFj9xbmWHrqMGzXX2pIVwVyiuyoG5S5oO
iJ0iVPbPstl8DZmzZI48Zxmro65SopY6KR8xGnnid73Clr5odXo0p+6EqeH260DYgzazgVqYYU4F
AtMJJJFzUhURHaJt/HfufouyVLtu4ffr7YXLWWMeEkTLjGDtWQcYrctm3RKmo7mq8rXAXysgO9Cz
e99PvXTlcH7nrHctTS4aR/MP8QwWg4ETNyc+asN7MIt20phXHLP9vO2oPDlEIk6YlMFJXASCZH3K
mZEj1lcyL/9jg/83jhBo/ij2qO047NtkRJsVkDLJnOj3R/xgfGUxxccxKdZ3l1wwcQLRVHPDQUhr
eMXIqs8o8FZt4cFXSk5uQVfSWECrIy1oevtZfNNTPkqvsT2Ytsmvm5CffOH7sAJRXC0n0If6GEiC
CvFR8WpjFs8fzpiEJ8rKspaonHFlcg9F7RFvzNixoHc7w6Kafk8SSw4AINyhJfH79P/CyQCk/poK
MUJgtG7Lj6E0jCgKFrDyjvwpaOPcObSfpt+rNGQpe27sKpqZMF7kMKlMEMovwDtX+7PlWMsKBh+D
iJJX3OyaXy5WfCTZO+Ul8Lx+G1KTU7MaZUztmD6T5V1x7Rwbr2grdNSmQzdUtHey2v8EoH/Z/L/s
wTpWNz6jGCC7ExxdvTZN2A0Vh3qsWKpNDPo7RaeOaTFlxRTYzq3PsJyGAEn9Ut0McXoP9UxhGy0z
7qlMOuSoG+8Z5B+FoQ5c/uLI+nL1mYBLRyQlgr03W1ej5fTnVbkfhdG30jOqnUG0BpzFagOLhqNA
sK3OZzSpR8tO/8NnFHdwFF78kjv9mDX1VqyzsCCyj2hOb4yT1l7WAfcBrwqPhjXpFzeFIkHsmt/x
GBaCDICci46ciaXFdFnbVySA2lxGnFx4JFW+/3cq5LpgUc00JX4CjzPEihjgwwYXAZxmAjxbcyDW
CfdpKAs7nd6Xzb+fXkaTXut4ybWOlWP0GMvMKQZXCLVqfPqX75JrwUGWpn0w1RxgVAei3MwWUlsg
FaOdYZq1EQJ2NL7jVdf+adkd/2r7rd1VBCA35m0lREyt/bewArKmhFmidY46ditTr9e3rYr6NBpa
vqe5LOuuHkPwCL/l3P5wk4iPMfydmW1S6rDgAHuiVlPu16GhKs+drtdrqQ71QByplHZUHYHbac6o
NU2NkIDNNvDTiLnMZdlLGhT4Jroi8VwrGqsCOxh3+CHyZbrJF0JHd9f12bI3Ri2nvLKz30pZ6Bhw
d2OAiZMOORWARiRVb13/riGOj/z7sVuHnRCAVutvjksdXTO+7ebn42YSqUz5c4qN+FMz+lhGBuzz
wx5MOeJCd1nKFzZboGbvOvrJnFT2VVQQj6jVI2LTcqsmnKbYTTUBs/YHHcwoXjAaBnyeTtzAAIzt
1o5Z/8flbBVfn2IZLexa/mXVeztOKSPR9IJO40LNMlc45FhGeKGZ1rnLiVyz0zIT3rpU8UyRIyuS
mEHfXiZ/EDXMmIbJca2pntJTNK88QWoyAqayqGctnETOkXJtdfpYh/uR4tKWdPZXP5XLZEsYUGIN
fbEB6IA6+grnNhZa4WTWgqsFP/+Lf6i+KOY/fKwGcSxIC9FhZAZPlbQ0fH4ThTWinBx3X4z2W7LI
UCrooynhhzVgB83jk6w9WbsPWHAhO9Q4S3dr0+UiBbHhtMOq7XA554NlSolnNQ7/VdRrBBhj334u
5nS1zvvXHMm5C8hHrZbXI1+mw+I80BsKROKRGBiPG5kLciAuBt9NcCX1MaalV7SAd+tiVZZm/s5u
oPOW1UMztOpKzZxFKfx77ZNmHDzRdL4RVIdY+u1jsDxP/RCOOE1cEVNwveVrizs3TMJ3JQPsLzx/
+vDmmjqeIg8mIfLTDTzmoN50IxEbtlG8hMgOJxmJu6dVeAHnxDft5ZzNEjdedTOLhjRZjiuCowei
UE9p1U8XPt74+chDV4MuqsVWmCvBOHOj6eJzWaMQzCiQgbF2UUYvDGyobnGImBo6XFb519Qs2B0e
B8HSI1fA4xrehUmsG26S7xjRlwb51kcmWp36PkeFU+1wVvxekOKiQMHdMOpjE7sAZ2pElbs0OKCx
x6izX2foPpH76YWwhRcxZfV2UfZ9rsct2HIjbY/K4HXBbrQyviZOdXZF7UDB48jsdzBQF3K+xk7h
siXoezWdrePJOPE3T8a8YcPRpZf/xkVSNZo3En84c0puUF6kjaxCCBkoARDO1/NidXCgW5YpJFbu
qCUwuwh2VT4xaYyDZK+8lmZCcnr8nQ66MKviUYu66NhZp8z7ztNA9CEdSf+yY3ztKO5VugbVkit/
Gq7ltT7pfh8RBYP8HbkExW31BTp7rnT1HBQyxV6zmNoGmIbGA+SP84+Z7VqaHejIKMIxqunLz4OU
7jfJAuKJfeYdbZ1jSzmoHreDpan79mBD3fAx7JW/Qnr2fRSH18VXwIFuBQ4x85BS1xQRbflwdpUN
vKhaqwmJhn50klt3WzWQzVXq2Slin8THwW+lcZejVm7tcBMhChh1gfZLJWDbapzSBvpMRdlveZsG
CvRJrtr6HCP6flsT2mzSj74qfQ+O7zeJ1nFoM/QZ2hzVysnWud4Qxkg9sn92aXyPeW8yHnPdnH+8
gob0gbq8DzoXdIt9Vi9qWXvdOsGo60GjsrS+oTFH0LU9vQiHbK1a+Fj4dNaUPw98h4r0n0RCSK4k
AeehfmSLzYm11+eb5B/3B7fHSeuBmJ5gWxi3fKOnu3LQXeKrlileiD29OfhgugXHI6IlNSdBITOu
RB/QPhZf4LuWOWj/r2b0hSOXGuLPOe83wMQCLE31h7VDdCbAgojJdxpZUNbi71dKR3pwZPWAMaId
BxTs6iyQMCEZa2jaXqJGP2IN/VJY+mW/QOswI7JGaDgxrZgpBVtBDgAvK/tRWXG3RtQnojvmiORc
Rq0zNw49IUHXppMUGD2BPjWt9gT2qvCXRKMrWqvZls1Bch1RPgF9EwDYXE9aAhPQNNs5CHJxB5jL
satlv0T3thlm/cQK3zT+YUSQLpMcDGXsan+Bg0OfWhq1C+Ziqov5JPX72QzsW1/yQ3TNU2e5nH81
qL+quV5lVRyaigPDESqtjA3viSTpv/rDJRLwaVFzwQWfS1ZcriYbeY2kRvwwgP+fwUXNjF4iRFBN
zu5wrDWEsp1PSBXHu7Ud7wZKDdGUqj+ZqQfPGiJGNZb06CRuw7XLcaK8CItlOS2L4pKjjQP3MqAp
ZJn/v0GUMm4Zb4VOiGidubUu+wmgS8hc5NlZgED6yeysYIrO/Otw7pQvx/Di5Dor7DOinUKOS7wd
84XI1sJGs9Ap3gRDiP426Su/Q7zqa/2d8cz5oDcRd8hM328W0M8NNb2tebUjoo3kvlK+EprmtCqf
pNQGgp/9MHWStZGGr8LYSVG166Uo+zMY3R+bqn1YZY+RMB1DNeTjAGeKb/PgJYtliQryFY5sMnHD
x+DGEpjpigw+zdzhe3bT8jqfJapdb6kzNEDfXUeS8iXGzdP9NUFqt5IkvLZqeCKtHbvm6yZPW1mg
8n5RA3DSxHZAywgZmW8Bi8o9o6mOWppIR9g6DRFvcUMqchuPpcs8Z3SKo00ZKpnN/OhxKVfMYA5r
te4SfaLxZGMCYiJ28fBdgMvEkIuBlQOXOdfHFuXJRJUcn5pFpjWKjLF9/zpsrbGi3w10g8v7KUpG
sO/pQzOfS1WjHgQsuSTSAA8pObgpgK+k4qTJLmdX1CX94Ju4fqNurpOx/nBznAgP73C6AeDbUSMC
RLR04ApOiUJvo4fiaq0D5B0bMaHn9jw/m8iOxkiCXDgPTT0AhyIurEoQyE73E1AOgAoc2ipYYWj8
NcMz8S3Ly5x2p7AfH8LBermJyMik3Vi5CqZMYodJlOEispd2yrCdINrIEneWSUuosVtTfIQqJaye
tArRdNWVeIlLvOgOTochlLmoaZWy0gy7hYRYswl1ZrgaNEIAxi+QrdOYPV0ezX9PJyOn3GcMBbwa
/BgcPSnyLoNRWelcqJfzH5XubSZw/cAcfdVnKSVz1zlBLKKEMrnhX8N74/qmsqYAxYizGfyRYTa2
9Qp2HIfZY3QH26+81fNupBgz5l7dbNfXtoGmhKX5ssJlAuQD8iEYsItAdYrjstY5cmGUH963o3yy
og7fSXMnhcz+mni1b1G/woDVwtBEnomnyfTf6dLjCGz6xcsyVBC0Lyj0v70Hv3ZDzUHPrr2MOmQs
hxJ9fiNsDTxB5za4Nk93Vg3K3vcRaxsDUvpGHbQ3o6JrU1qWoUzXp6GvGYwQaykm5khPdAFW3RXB
U7seRpMS3QcuhAu25GwZDSrJ0UGLLC/QRibJXYWeBPrnBXH7bTUSQHsJ6nrc1jL1j8nfAOr+OGpj
ITAaTqr4DGyqhOSo0Smw+67Cddp+rzjePC9DKiTpFIJk1sjf7HwV+kqtPRQ4jrGa7yR5hzT5gqiA
J2kztjl/S66oZ5C8RC9oBReqKlhz2CNZTaHtEKarVASnkraoUWwHztWsG2HWWiNUzYHnNP+JwtoA
d8GH/00cTIMP0XoefAKRfyX77m8TpFoyr/v8FjZWa2NkWUk7SNJJHVgDShvmjDxSTF/KKEImeXp8
DFjelM25SC2YOiigIcpmoPYefLJEkweVHrikPHfbwh/I2ON2ybF4g4qfs5Luq5XWgyWMbp27UZ6J
GEr5EEg0854L56PAXRzGttXebu6EHW9v0ETxyIiBMIXX1Tr+yW+YksHngPGIxQp5mvrKiSFL67Le
2zaX2fLHdtiUWOpxjxa7ffK8FJI3TDPxixIIU3wSbOhC51k1LSmySYqz4uFfduBPS8XEy/9CGbsL
UDKB90lk2bIdLHgeP5ielXwegnA4ln8XV4VU5Wt73mTgtWoJl3SOlseQEzNJiFgJsItNQ3xNa0ie
gNHsEZqLKh7WQI/4abeeSgFD+Oeqr1WyCjeYnK5LJgsJSZRkhkXrA1O/wD1WZlQ+Cpax8KRkax6d
+6LelMYiJtfaqpO+qH7u3aPveg0U4/43CWO50Ft5/A7d9QohggESxMrAjyiJLurQ4oW1/26SlNu3
Ek9BKnmvJOD2j7P9FuA7WbHe8BjP4U6gDth9Fs/yO0WPglwS3b+4fG35afCUdqoP+eKk3j143s/Z
94wZTxR9chZ4MlvGWU3r2nqOliY+MPW21ZKfwCmWCKHozNuMMHvnXY7ZLI0E6Mwgw12o67LNw31e
UyZ0EY+Oid7NPTNvdV38tFnxth6X+xuDvfbSV/3CBGWMmWaDOBr5lJToq4Q/c1uvt0w8BjD3twpi
fviUkVr4r1A70Ypau7HzuwlEqgfKZj7IE+BGfeFXhqYsiIvWscjqhGQj+rPdD+U9ah/tTxe9bFEV
NMnaKGx/Ky06axhHeE3h3OxM+XPSnN+CFdE/B3JzuqZJSiXeHhsfpUecOuKFkHN4w04rSJNYc1Cl
JSa17jNwpjRDZMOTek+Nwpfbaes6RvjJM2Fp7VQha3UkIoJMVgOAHC82gMpk9Q4aQ7JA7OQN3yP3
BaVoOIDrAHTjqiHlo5QzyOEzHgP5cfYmTuhEi+/yaWfkmD6ArBFzOCWVwGhCcWOH5pggLh/c5QJV
C9SNlzWbkdJclPmX9huk8377gk44Mku/v9/AC7HCo2FYWFWYy37IR4EQN1AOLyTdEaILHF2CWJOD
xNwmufRt6U1yRYlvTm8Fbn6sMCeV7LoJd2a2TZqoRapr25k0dHUx7c94OtuvuRk5jRBKQ2KOHcHy
VAI+uRu7iyXYWrJqH4W9jBF3EvjQ9hlTxQEF57tlzLNYgz19R3ZaiWmwyxI7NmmHg6F5UldQD+oo
5A7NMrBuJJSnrc+0KZERd5XL17TJvnQKzIuEGDraYDWI7f+WKRDI4T9NcyDz/tZrg4GcpCpEImSZ
oytG5QfjPK4CFr0Yq1cKxIl+uy4NDw/1zU+9fRhOadkhgsKBdtsEwt/q3a0yaXMCuK6XUr6OFNP7
oF0/20X1ESk/VUubXQctNVrBSz93oh/FtL/zWljtWLi2LeT0M4itWTV7LU03DLYesb39yaUKKBo0
ewKqCUxf5bz6LNM9crXbPtaVME2Rk+Opkn8XBmL8fY8aKpJu0RDYFXdlZixHpBAJDCnJZyGd9slf
HUk3+CRGAg5fl9w1439fSwyLLcRBe+iHTa9w0NDU4shAcP2WfpHFjbxlbYvzADUjmQ1k+8BcQz1S
Qdk+cUUUjChJXwLGYwha7hdZjQ1zP1CVsbk9NnGg70RQKt0plkuB5Xg6eiAbumgPNpSkvh9kJyP4
XtOuOiU0m0B1PZCxJQeA65ufT4EcxoUwE090Qx4yDM6wNl23NMf2vg0eVE+ZZ1bQuKcnejQW8K09
JcVC7E5URwgoIWHoakdrUUKDgIQ8Qnn+8fnB+g/VkpOEY4gNTJsVqQTVUd4EggAlLOoFL2hwP5Po
bv8r78cPQ2IQkJm+4P/ay/1H0mRi+8Pw2jJJbVcFxOYnjqwd4bZzh5wdL3LuDvmRuvbC/kwdslia
SQUkvVknF8s7i5MG/4MfaPfGxfmF3k9OUUttGI59FDu/G+d1WemLjGaqW1lD0SWCo8tc7Bvr+LDH
EHtAu4OIc+Nk9U5G3tNJ6es/GJM/1ifolHTndQD5EPa7pkGtAwL2m9zWZPcR5dHbn5QW7d1+yfi2
fjT+DrvHvxVxaGq5hneMfFMS4zDaAB1LEetJIRkngF93pG8h9hlIxUDsAGTdVMT85LIMNNY/7VTR
Yk4crJ1MVeK5FhaFXjVuLb6xcIKuUscQeWSXJNsnCbaaKDlcYrrMDxWUbOAQ/Nx+sWwPNHvh6VYw
O7wkif/x6mZBphyzoy6UG974GK8OPmot9DvWZMOdCnL6HeeEbgDvRL+hHBWKbsKHHZwMj0jVzg2U
HDzaTV+gAWeD/UUsGss8+yOdVFW4sOo1klSTCQxxDRyQ/tNwGRGMdPPPUvyLtGGNMS97NGprzaOB
MKHYjdp4IPL+bFomld8EoTSN+gHJTwZADOC9BPesmEtqzEdVSHdca7EyM7V1jiyrKUSKcXFMqTNc
k31p/C0NiXilqy9pMG++uhxw8cuJJ19gXFhBTiELoG2rt0Lj4MYO5tbVEGOxPg+RZ3xi8wOU6kWj
J6L4QLw8v9A8VPMFXj1sLLmHwvhtYHw5LRbOuZqO3CHEBcJ1IVdmB88Zgw//s9LqhFrr5Lwsy6kP
GycSlx6MVET9j/HNwAgSAAgyI3BMptscaBh2FfcWbQ99iSKzAYFi2/yxaNysJ5VXPXuY1nI87qUG
OL5wqF3IV+1pfljVuFBpOvO/dgv9KBBTzoFkT+Ji1jGZORexOhaexQv+/mzVYzGfh+3v4ccuOn84
z1HxCWaGXodGao6cJZR9I/G9vfIIwo7hp+JxEdWXhscAVL5m/20ofHkRXOKXSSJPiYLSqYZTrU8H
3uZ0VqU+b8CW12PZki3ewr/8Z7V2jC+V+7L3lNfRk3VQX2aB7j1u5UPz+lDUG0Zw6bpX3+fJSEWZ
7d17nCPyrLzbALXuDNaUQNWgwQjBh0zv7wdMyz2nabNglolwMKNOegiPq2fpYqSrsBO0omwbXroy
K2vnAOXr2zKf1zB6FO006+nqTPJQf2+pwNp8Zuqa19hNRtOrpPoECUDATpr48EgGcVY5pyIpLQ/X
cgHx3wR/rQBocdecQeQHNnVO/GTvzTh0BfqCHj5etwX7BHeCpu3GjZ4zaGrE76AYwsFinpxfQ+A5
NEa8PuMa3LqUMKCbuDw7omT5tH2plUZylGvwfjLse8fCdZ1HsGbgJgt7lg68dbTtPjf8F1c/gg4a
zHWZ5UkqeB4IZH8slLbvYsnFzmFnq9z8bLLSjOzdhlU1RKZkXSTO9AFwloQX9+cjv/qlMi1FMbYl
ebpGSAiQK4utYEFJxsgm9CeIOwEPTkxkcB4dVFG3hzq136b6e82hD9lymXSRzA44V5OMIYbszlTD
uukUoJKoKwiskh4OMQa7vjcmuKrjkgxAYoFNAU0IyYXkkUfBemooOzusIdt9131PwWlDlxTMOL3V
v54kx/tfbcK1CnvoRfs74gdGIEHfBAmU+BUj3uVIdbgRfGmUACIQkVszVnMLq2Miq86Fk0W5V6OX
IE3R76NkoDw0NXA8xns+DOZyxuuUfLG+hLHVCScGFvn6nxN9gFXBuNH9q3Kl0b8ys8GAbeo/Xo7s
bj2kwi6TjldrZa55+ensENpmTDSyIId0FpsM14alpaqy1vPKly5lLixuTvzYxJq+lVd6wwAJ7MBc
Y/PgjIc/CXVxQiLhI5O8M7kD6PY06A8iGrXuS6hbEBnF2tD0BEBSezVzMubBsU6Zc9/L/ujOLV0c
O3v0m5fHZYEX8+CeroqH8CnVzy58KCdSLqi6Hkw6rXeAYaQz31QZr/DgoNYZJoQjiHRSlSk6ZoFq
Mib6iPGN+ql/b0qcdCKzu78g+3DKpASig8rjqSf0kxZ68Hx5P/DTASbbrmf2sHBzLTdI+PtX5aPA
ex9YL94AtYw6FZyOVxZsRLH2dMV5N3LPGSfkNBwvTitdbiIUWZUaDeJNr0fQQ1ut45DTAoCwJSs/
k8wG9yb7yAT9mLrrI/0jJZeUE/mmS5O/EdudZbgxvFt58XhD++rYVkPNPV5s+orSKLSiqrgqelWy
KEovLBdepvioCIMXw4BojiLQIEiTixnRHADpPdU8nmOYqyIwceyxMTH44IPh8k3ML/0G9SM4liAM
7ir8tgDpVvxobohU5h+NBDKv8/jQI0Wldl180uEWq7uPAx50YfecUFTqzSrmp4ihpu8QqbtCuKze
dxpGuove87usZUIDKELwv4ZHDRDdik5FgU4714W5QM9BWyKDCAUPFXa8D5nS8fMDxpWYlMZVL0WJ
iZfV3qtcGzTQvMYQE1CmUFib0x8Tuimm+aen3uTcdRPJ+ydbH83Bws7aCRCqWShnAsMCYOjEEQQE
Y7s4L/6Y9MdWajZW11wwCrfo37FCmgoxnqnjoDVIUVfwQJaBV8/zmw6AOgNuOJpCfetOVtGpsOGX
05Ao+QGmTUDQ1A5AQq1WiE3ZliSz+VSXBTwcdh0A2++9rj6LkABrP/8wua6bu7m4TIyPYJm9nMYq
Cd5Kw6Jq9a+n87mByq6uDoGrUtWd0fMs/iX7kfaHHpOkbVKUVPJeyNdzr8oif8Soeef1FpPbFyqX
oTdPOoVN7JscoqDAlvoeabBF7JDVRLmQNUwiUsoKIGi96jszCwL86APiVhhnv46e3gsOguX+wI59
Zwg0jkpl188OkZT2wpkh+gihARQm/mfBJlrrKEdKixX3JskgjCkc/TY5dwFoKJ2mWZTPIxr4Sdti
Sech3pLjLEAF+/5jYCdBMPGjaEAufOP3RnaCvRD6O4aRO7IAh01zTBo3Dp6pp88kC67z4+9+SCc/
+GJgpAF+OZBiOM/EGs12EZe7Z1yxEz8TWQmhBCm/UjZxeIm8YuyoOeAmVJxT3Dg53ZK6pwWCcNCW
Jvq+N8MrzspaPgQzfyZKh8TVp00WcuRtkqIOHT+Iyg3859ygitzOq3s6DhHUyNSbZzLgeccNqIYF
5TRlPeEpV5nBYRFNUyPFXNTX2esJWWUod7rC0s+iYQXIjD4h3xtVYmUQHgTJez5n7ZpSGeUcMvz0
g7oUjoJWxC+a3GJX8tbUjUwrfUj2eQVMGDXN5uqESBxyDL2xERaOIqgseANBiMye3uupbAkO0+u3
+i/3xCvaglv8RMXCP/m2XSteZGs6hEQX2CwIpe8fOA2kAwIQiNb4KhZLfU/Hu6tqsntSryOTPs9X
ovYG+DkjycTNYLsLNk3WBRIY6VMJ5CQyW33+7z92APRLg0Gm2tFm7mFcwkD9LqEN5dzd1A79zN75
wOHEsQOoIwOAesHHRaR4BvlCZKPnu/OcGJpj81D/pkJ/DF9QDaqgEGFoNTcbj67feVrAVzQHLwxt
Pgb7WusE/0/hiTWzmhyig6lALdDt3jSb/FAny3OXA8kFxPkkYoViW5eJsBxDQNwJjRGJMOy6xg8H
lvVJM+dwJhDQ8VjzviJWhC5yNLNQK1/eIYldrNLQtwLncGjSDCy7bw6Q/Hje/QPWGc4FaaiX+9RT
QURGMenXhRGzSxTiRb7AJV7Rk2HBR+bFlNLy4Bsp+PkV9W9pxTDE9f8wksX+MIEfc/ZeSidF63mu
IiqEgKGxY+v1ZxsGPl9Om9XPleJZf+xwb65VONmStvVE1DEehcq2TlE2aSh9LErLFWzsbwQ983s5
N4+EV5B9c3PPpEwLguHFRaFeP7jAI7w6a5PZ6l/LiRcLk5UzWBN69be9oFJOk1QicHCdiRAO73rp
hXBpc+HFnIBraQiLeEVx77SCuRtAsPsdxRU8T+jrvNY0PLclCzn3mAJt3gdxQWP5ZI42Ktwj/TaW
kbCtyv4yDeEjooq3clnoGydyNGqy6PewR+IREutM/pzLcIS4Onbogr0QO33JPQ1fwacpKs9eCjI5
s3MgLgYZRK8GUs2Mw98KRG6tuzQWMbEYarb3iX8oTn66ppSLs0gVVpJxEptQhMSvmK+y/ng6DslK
yiLn8vayvaoPtuBfzjvCqaLjYb/JPZstJlt0kEV/9lM9OeHGQdoQN8iCFK6MDJlo4dFzCfONQCRv
LwzFtac/xI3/09BhBBRscRDA7rUU3I+ImlsYglMj7GGGIyY/WeVrZid9U0MGR/5sR/mv1A1inLpV
/1u74ZZucmvf5Cy1blmi4LMDGnX8FsPoM8fW9yWBYAgDZOUqftbfT/IP8jSP66Rjsmlb76ZctFhY
a2xqCNJoSEirH+imolVVzjf2t7XYNmgDyBkSeU7+wU4v/cl5qv/3tIylns0vjhy3K0zV6R+Jtkhn
8fOjcp22oyvsAO40IXpjCCnrSQvm6dS7G7v+oO1T9454U9SSMjVL2iyd1WAuBEqLL5rKrHVHFyCb
mkKbXBPrqIgKizcTRqp1uarJtK+8dIP1JOzwezyrikNKdTBDofcgwwrT366K15vV3UiixIlgnDn4
blV5I8tP4z2cyDP4fO0SM1ZBTxJBRE0GDO/qnZJUtM/iLMkX+o5wJFK/vqeFd0y8LvVj+tJ8KNkR
8TnyUwef3NWgGgmZhTZql/R6jWZkZWiUYEOHRhrRj4/YLQWJW1/9Tso2tai/gZNbajpZ0PIC+QnY
vyO6Wg0Vh5lkCcLsVphva4hPJ6za4MIXInbdU4jdsEsKmDe7OV8ar2qhUwjGeoAKmzn9DQjkGg1G
638zFqx005YTDsCU4PikIaQQvG1SY9LTK4D7Nmkj8ZISLFTHedOoYkHpCGeq/k12faIuhK4tLVcA
Tt23XDxPIxiXtHPeuFxYYKRpCt2ZE1sqUJO+BdEu4aC7TaLyESaJKsDI+fXNyeIS84yfbgLfd2g4
J6RDia+RKIuv7nRTNiptUwhPVNCALZJTXeiE0qflHZiDwSPwzxWPyId/jrtVzuAUBJM9sSdGdGA8
6o51HSQNUujHlG0QXCsTv9y5MgYMHpKK9W7LK3c9sk5tWFR6Olo0Zv/lt8h4eX/tlpLD/IlOFvmC
sOjAgKt5356MykCsqh/65mOLjrGK9j+j9wRDPh2Wpu6X/7ctBfiKFM7ySN6rS7rTj8rl9xP9ssMw
kiohzRUakgolPtKN1NjPejqWrXXWJXBfXu6BP778gvf9yO87nYUMaEQhJ/XLZR9j6HsF1b1xi/Ut
oQQxonPWiuG7WEFR9Ciw21NYwOsnsTDeU+jXUCkrUiB+eMEEh8Gc4EneX5g0pKT7i2HBwCvCs7q2
fbijXcC3ykMR1Gxp1kk3Rf2EXKlDUTknw+vsj35VIwmgqCB0xvilFHvDUijB3rZXTOfYQoB0IAik
1Ea8oNf5AhOTvf4PM0PktWvXykuoG7bcEAf+M9/ojnquemNtxvzd3fa+usq08U/n6Qw5M+FZT7BQ
Q3m38aGi8qFKYAdbX5abAkqJ7qfaGGwnYL/Cl5U2mXJM8OQ1oKWVVgLvw7xM8unPlm4vpCOAWoDt
UAOHdyYP/3T18/OaK8u24daQUnfY8Eck7JvYRtKcVnXwXRqXQ1LxWxse9Ut67oo0ZHs2xlJjj9vV
Fm75iDMtPD0YJLIGnJ95e99NML/wxXnfwb6OhffM8zESRcLPGZBE7TjTPqlnsbe4luvHmMpoAVzd
wNNoVLxxa8txnu+BWCzNPcY1FXCYWtvX+EiBE+C7JNYCKYRFgYlpFQZPqrIoyk20R5NI/WG4dFM7
1Txs3FdsihlGM74mtcSyme7uhicV+sC5LjYh37PuWOMGstxu++4Frh3qZMzAMxFRzZxia0RB0c87
ylSsVQpaSXPQXQlZDxPNt2sdXcPLwlVr+RFxaCCVPX0+wpwVV2m7cJLfROC9IDpF5EpvbJEak6JW
aVfpg+loXXYRbvZYO+iA6MZvKyvAPx7vMNDhPZhk6vAJWiTEdtbFSqfNluqPCj6YN8qqUrYum6K6
+Di+kxxqlpVUkY8XMiED9CLmbAW7BlXSQUqdb8S5gmlKzmoRh793UuGClxVdR3gAnqTu2ftCgYi7
96J0v+qV2L8ZhomzzcCErJT/f0yr3WfQrJL/N9x+SiggUhCINJeozUZ3dM6gvljxvlt8DuF7uxTz
MsreRxzf6L4pllfaYImHVjpuLxDvGJ/98qpex/W+k6Jk8Lnu/ZpTUU+uluadb/VY4RotklgsY9Wu
PCmRi3PcT/PM5OqdSELvYxIkvKEuY8Xvdt6O51HcnnFf6HTBSB9QGceM1/7Kb+J81qgRVcVC+PXY
wH1yOd9WCwPPD2k3fYEjfaNQsmDX+BD/WqpbFsoOplWSgeblvoKrv8cvbqnuF8TM81CrZQr5idBx
ivQFVujyYhjCSgzD1Q6o+fLZ6OD0DlsmFQH3J6nfml5flMljySkKqb8SqqBgxC1eVpG0qIcm6v9y
bCTkcakF43Fu+Gvky0RRhbcMaLFLKHEyBWap0uqMGeGb6WrtTv7OOCqjiee6CjFHWJDk6JJ5JO+0
D+13Yqj98yFdqWlCgkuAgiaw5Jg6kN8QBwFHDn4RKewRBHjw8Cm6zsBQ7w6+y2sIKT3mTZ2sqrz5
YtWHVJtJ/lxq+Q7FWV8GCRG7qJLWCBJWZXKNY2Fpm5Pifab28caGsYC04ij75mHbf/fHTW5b/qRW
B3jkqnVCXqRM5JkGEIkvG3ZDwn2WJda+A26Yfg/aFNFnAcWTiJtL/d+3B2edl0n1cfCWc0Td1Hzp
thy/4RlI5ha0ICBVT9T4TrcSsDtY/B7ED5PzYsJKeGcDV0RVX2E/kwzZu/SW4eMuXzEhyVNAspjD
x5/DSoSr8UqBvHK7Sm3uvyGs6MaKwTB5KA+CtBtnaJ7pnEbtf2N/NEbs4PUIg6wxhelPAbUAQieH
N3G43cVHOMQ1K0rKWDj04YpQb8MZCfBTHTuEqqb44BUg6fhI++OIjGQcthhuTIlOtSCyCXljRiKb
E4c0XTtlFzvF8wgyTCJoLoVkz3kul4PTNm3B5w+wmXRoJ5DrNb3wZWOaeVRF6QGlqqqc22RVvuwq
z8QC+TmjeQt7qb9gZ4gyJTW3NzGSNXCaG3Ueh0l2kjtwqeosDNgReBgJYni71rcfN6h5kMaim0GQ
VQLudyI41hXUM31WQ525I03tOSUxh0TVgU9gygiaz0e/NzKPvBb8DpL43XwLmjEAPtzKuKIRlblf
F9d4K8MhZmUaWQvIrtrFD4TFPABMvKENbdfUQoK0Zr4F0LgPSwkjcrBSRkRCMRmNGjjN/gcrrMHY
/oRXtiVpn0XE9nDjEFRGza35PzReg/JLlmMFg13J38h1yOrZ1fO/Vna+EFI89IuXkGtBi9Lt7qZf
8KdFqAete29s+llIaQwpdNazJwLv7NVgU0KL97KaTHLHY3ej8khxHaUH4udip1+Y1dBxhxzjOo51
aX7i5KO9PKEXzpwezBB44baV4YjVOt4oykGn2uTbDz7tPrhlhiJJBv/j3SX0R+J+NzU5RVbt0Ac7
Y9UREFs6PVrMRoL5SzQMtAZdh1ONGO8HfNMX8R1H9crPKtqooeshn6VsH+bAukzTVtoMsS4kF/+T
j4uRB2ZyMYbknLQKTnl2hJCjymtHvT5DhVB+0L0rLWWtY657j2zpQ3r/6Mq6tGwGPd2tsSgUzYwz
GNlTXGr44pdQGiE/k9IO+YhMZLoYLhoEkqvNB5VWqOSJsES9OPDQywzjQWfbHkauJ4s3J4vTnrJ/
8WxHgV18sFFybWjjFb/sYZXUd+kKJRFVVFRjg7wCFMK1utaRNxR2MVqgrA8nmsFjb7CjUPlAv4Yp
Gskhq8qRLw/ZyW2Zuz+g2oTzlGICIUxXA9exhNpS8AA/WzRBMGkjcwP6ZDy7asYERU/pN8leC6P7
WVtu+tkUk0c2fgScz8HXAzszpXuAT+E7oPGhoQi3d8MhUF+dzA4Tbm78eygPsfoGuLEpwXdA4mFN
4jBfG6LNf2yNRzsMcPpUrWtQWcS7WU3KmZ+aNGF9UL1rzgzzR/Ndd5OzLF7cVS3BaWbkCtB2yF/b
H+CL1hSBqK+dc0Z8L8D8nutSNbdXtvw0AT87zuoXZw2/Ub4d9Ws9WUXFgzgRq8zVVePTNr4wIVNU
1XRdiDK6XvR+j3KrLqIC2yhwbdYt2MeIPx8oUqcg5s3aPYhW6V4IHidUMVOWKN6mSUhHkhuTCMZ1
SNSyopma/B589BVqZ1rb1INnaKEFuBTdvgBZWAODgMF8j/PimdeMpaPzFqNZH8WqH84DSgskyNfY
dNmRa3P/9o+JXLuQBKpUIFmOoayjTgsGI4mZjPSoUHJ9iHSqyO6NUTmmkf8MgF2RguA4LLsiZe4G
sVwWuOgWzY03+i5h484faYFBlNaqyuQBZ4Otni7C574/2MVDwsXboZgdFOnXWRJkByBrEq9Csqzy
2ZVjHYvMyJO5adqX1XAEnDrFxhDDjHwBSuKVxkk20jaSWtKKcb9ItMU3P80ruJypsWLxwgxLkUM1
U0SodqUXH0nfin32PHgGu7VQFO21T+3XKPYJf3eWIq6eyBKsZbLE1kRDPm6vexHU7Lc+yWSryRDU
6au4l9vOgqeJOtbUTSErHYHC5BaX7NcscSWg4+dEJYEV5fXeWk0B7imJDCQ/Mue5Fwd2jo87XVUg
QDQoTxf0Orj6OWilvR7l7cS3nB85Za+dPKHpK9l/zGAltYyo869cHAXQwTTF2MFur6MHMsqMEfEz
OxZM5pFZtcEm7igy+WKNYjWrgho/KjaCCXa1pw97JE2xOPVm1qTER+mQx5IvqpMdOd4ohSsj0oOj
cMEM0QiScgnfAPKWWxsSeA9liWigpfmOzAi/dJfk8oSkbjsdgsYiVe+zb4R67ueukOsyROean3MY
jGviKZgGdUYHbZ8bQ2kEn6SYkrskwVwJYPhRj4BKRXPBlWf3kxW+Z5V/c5V9VvpR4u3uv5deqRyJ
EkS6A+sbl4RkaEh1zFI9LOe4vGnn1Qs+pgUFe/fsA06dOoK3BWrg1TDl30KzNnivoC43G8AKz5x8
qHbwQsLA+a6vFj8IT+NxXkODcIvqqeWLcKDtsxA7yvAyLuSoyCSq64d5JEYKt91bbXy8D7iU8sSG
vsF/US8t7muwvBlpGyawiHQ4PAHwY0vFF19yP680rHphig10KHxFiJZ9rKE3h3ZHi2N85lk2xiYz
CXX49D60ELTyHWvpnVsHHeQflshc2J4aGK12PjbCFKQp6NruTGnGC3MsdxG4OzZx6g2Z5HczbGnn
dx8uy0ctWUQ6Mz6Kvs2iBWkOyaa3rXyjw2MhKtBCnKUKcvZ2uPYZ1VeatfUxoMCL16TUR6MRQnov
mDC4syQatCSpuHYrlDlya8a4kvNEcIou5t1NIc2VeE0S7EFFGts/EKTNvyN+NLhimX8Jo1IRACVO
8ClgTC+aGVWd50CxDkg+ppCNYnL5jv/UgO/QvTbzk/azgLhPW1sAKf8oeOO/jV18JplanKN3F3af
kADm0v59mM8Cek3IIGM2hKy6TsaqrEVu2Of20H4psmHk8OVSWCUVv6YLjyP80PqUiru4JZOVUx4N
eV9jnz6J9fzsqa35xhzh9WKh7UzAtFOUHz9RenXy0smE9y1waL44WrEUbiTGd0QUkSS2QsROqm0w
hg7S8VW7/AIEXqhxg7kLtJtvzUhQeUY62jvDgxM6byJ2GNoe3wGBxeeyIPiWBPdKbJSTzoum1mN0
Fh7FBmWD5Ecgd62rQlYey7gkGL+PbylnJ+tnbwsW4QvS/ssv9kq3ARzdGk79MmUzGs6DFk+XRBxK
Ew1+21j4rRfGFbPJNQu6BXy8jjXl6AboR3J3BuqRiD5JnRCn4Zvnwuu5vlTCtHDcvXBFiOdU8HHv
9Cm6RHTFJaS9OA4RjBPwtfWtob/QJEdyQ6B+ssj6l/sqS/LVjLUhgKqsgzUPEuQqIksB+xuNi/lC
kdMsv65KOxt+QX/brVxCJ8eNF5C7rqD8MgozNOro+RuG/4VjZRnzw1hTxrigu0Hq8nIzhp6grXiB
YAbh262gVleVMRTjUBO7dPUK9NN8ef9qrp7BkCqlQPq2q6a9ixgfHXD5HIRxRsE9vXagBqBE1l8v
1pbXzYxfGS1aMPgs0qNF17LhheY7mB/mWU2Bmo+0H2o4uKU5BeMN3GbLjK2gxBrfGPimRzFDQqIm
YW8r2y7O7QtAaghduKi/mnUXhF4zqtOsIoRTMI3hb2yM9quYF9adAQfrpOzbJ4WcGOoW1AokAcoV
5gmtcYw0JiSYOsmN8untL8zgZ+X37qtD9C0w2AwVsKbDPxURaufqsdurltulsazTzqtIh3OAK9E7
l31/8wGsABH2+gOX7Ob05XbgSasJN0XYW9iEGOb+rhOQRpRLenWYoKYFp1bnG5Opp0TJ82u7IVVJ
xMyyhZmM01Qt713wRp00k7KNjhR6oyudnqz/ym2Qwq2zQ+uwuHw8usXAqkH53fSEai5+EBuOZqms
OBIOvuUeHhM8m65Uhosh3m81PNcCEdV311FsecP2Koe8IvuhRZUjUsi/ssNQS0576ffMRvkzDf5b
63jLD3d9mZ9o2elgrWXANqwUyMI0BUptNvRu0rM5LyFGkthqlsbe0/sVbrvQry4kz/Nb1M9t2uOy
3b/5CpqMf6pbPWcdVgPzAF1788MHdojBqv5xBBsrmF6rfRTsd3UM/+3vSXfRT1RM2ffGR6MT85Nr
NaDtAjL6H1x2B3ph1Xd6ZCIFrKznTV7Kj3tIPG71iDHtte3zR/BM4XetS6ZaGQG+TlTkNh4PTWim
jKsU4Au/Y0MJNrp3wfRIQhwmhMeavf5Pk8HWvDj2JgNrajTskpx1AhWkMSeaBD5Ez5SjrhGnrYI/
tvQ6dbIuvjzy2SdGkx/18RLNK662CCJsPox4knv1ALr0mPznUZSenYw5YS+yihu95EbW6UUnN0eY
c2H7ggvnuKPHec429+gRxb2RXekzTNbtBh8116JdlXmX7AcGQlLLK2cyrpZRgYNSMgYQtsgdIPud
fVcELtyiT1Wmh94R39ZvF3bPUlrApwr+RvW/rNiVf9JlQmDlzJae/zCP6SX41MKpbBPTg0u33ZkF
j27OtPU8VHy4dlWw+OEysWj6rSWsbIgh0q5/hDf4Q/4dYkjTf2DQhEN5W4WaIaxJZF+KUHD5Xa/f
38sxCzxCtD8N+O3zrRc+VGnuFfUtQc/S5kYWJuksadJtZF/Kya+sf2pmnzquScadralrqgdPFDUU
ppYn57AnmxkDWmhEMXyxhEMSS4TmrVo6guh+024WtGvRJFqKe+eJWxUkK54/dT82U1QGOLM1b4zJ
PhlX2+m1zeVKg/e7nnNpgiZn/oPND6gYqB8w5vIWjN2VLg0KRp1+CTBWixL3LCTGa4KNky6SEG1w
wmiqt6lz3MXT34c5g2PTeg+Df1g/D00ZcvI8nH3jr8WHErFwdOClKVkHn/x7g608kEMlsTviLfYD
5tZyhw5W9W5yoZsr7MCgxFvq20VYqVlO2HVUzxFPpH0NwAghDMelLD1REdHnObFFr7yIxM8rp15a
w2/APM7Pf1gyWMfaQFOcg2F29jJFd7fmn8JtLMUs7WlPXP4lf10uuVGmmhnqEHacKGmd8JCoZaMl
baOSFNDMXDfjCm/NlMCWGlcl4BFPs4vg2DOIelQZW/qpA38GmyyqJxBo5MKxpeKNwLLt1V0veC27
rrQ4lA8lIc0m/zpOv5HyoilrjwPbh5B6KIRStDIxv2/9KBUmohQLTTKerwjz8cRYa0dZpHqJYySk
2IddTMzurHhIpab8i7Hq/XGLY1G1p69T4GesR27i/WkyU86+DKoW9eTxxHlGglVYCs+RF8G0pZ+3
Zg67RPFN9Ic5bPIfwWvQ07ySApr+nrn3anqNA5dk9gLwVJd/wYKJv/O427itOSlnWPFF8nQZgqfm
v7bowCMhXro1CDZinHVoBaqEQn6xRwMrXOhn4LvdKQlIw24b/1yDZgPM5GUBEeOQIKpT+ILOvkX8
afE/IOvVbMvzlktvs+KFOyQ3QtJZtepl5Qx7yZye/T0QXyz9CYPW7UUyfSf9mqm9UuRxUuX7x8SD
18DtI4Khzc6ejg0QQVKtIufA5JF7rjrklR/YsgTJMy6qkQWlRMsnPeGmc7oKAxfLI6TnvaTAluNF
9nLPuMPSY44HKPU0r1gwN1oDtqPl+C8ZkIPJ5IxQoRuN5Hzb0nk7chmITp9d7hVF3+Ql03ExK1S0
n9soU3fRlxBScre7eUhC3/9VkeP+QAppyhTFtGaNtOsb9ezqYRt1tZ9Y21RaPU9SJy5Kzxdj+kJ8
xHxw/9lHAB3kGuQrKsDuj+twwpdUfIRkeHxUTMijJwJNg1DOSdhIyojr3OoGpWN0LDjWklfVZHzE
TkN1Fok0c7H8+S3WdoxekQ+FDhbd/ScicJ8efXrKzvGug2T+6oHsaLAibI0gS42mxP52uk4QoBFK
+4bMB4/HBbounLPGUOvBDxFUs2ADcAd86cadnxwUbzMuTRh3Ehfl71P3xUisU9MbWkoHpfwr3BFJ
ViykBmoA1vsw05CUteEf9uGx/HexAuxWI2/rvphO6MtXG93YMjJztanHMY/83HbL9J8byX1S0G2A
LIVSBxSR7Mes2jfnekD5+L1yNV/PxsVfuVkp3O3sw6jppqGAF7w6F83PoubaGNIpqgkYvRbBWEta
sMyVvsUjryyM84IsR9x60l19ibBPFZlar7K4Rxqy6DC2oC+0BaTnBNw85ifybDOBiDnmUFwMadTp
0owHYTtAOQ4/8B9ywZgHeeg3jJP7LAZE0IQP6PVdeevlTwj/+/Bx46lJjqjGaWQg54Y0bCczmXqM
aMgC7jinbPuX9wWWWP0jNKAv2+7ji+zPVn0nUqG2594O7XmzbOnm5VcKpduSlfZRnLcbrkmY+Qki
5AydrPjfmc9UBdwQK8bj9Siy84ST8S3oNcoik76iT9tY2wIKeW2xFz370KDD4+OyOnQwP1chIpBp
Ed0oG5TQcIti+j1gmhO741bHU1ULEtW7trteL2U9rKAJ2sDhQ5a246uWSHAAlzRS6wQWO1E9/Wu1
CXKX7OqiaZg+hk0Htiz68s5B34ke+IUL0ZXfbAjLcGQfOamaKWJRtMO+rUM3lJySxD4bPktT3PrV
8n8DfsSpM2b/e8ItM7EKxJB0tvMgIjL6ZOuyCS8DO0vSwuapOXOZaP96zilYez0aJutuc4lVmK9R
MYcswHmkw7OwhdQDnNzDAKZOb//dY+3QJJY757GQAmvbGyvFB/abzhlnO462Ie+BvpiRz9xHeDVH
nLOzhWHEjAqYBArkrNpU7Qk9BL3DWLGjgD1ZyHD9l9psZ0eIYJjkkSOhBwN0/3OsbvkRFZlngGZ2
3ulHxI9C9G7jVNXs0yRJf2eQNnSNl+krxrHvdtW/4hyEeTfVz6NgpxEfZhwAKrrp+kryn33VS2qq
/nHAkR7qCHqS0indZbUvxv308tEFd1guWe3eeZ2NMLqYPRHKmPnpdn8YXIf1Kk0GOhf68d8OsR/A
iYlJlEbd4nsy7LRFMcm9qQY2QAYy5FGoLP2roqbWxdutrdqH88JhUNAHQQ5j2rj1TrFGLJYCk6F2
kUcVfL5+0qLsKTzslpHpd8+A8ksZJJAugmvJo89tnEn6GBjXiL3LOZzXwpgi7BMVCbEo9h2PPqpU
X8+ULgRPr8qRtySY8oUuutM4Eqk4lx927Ili3xmu88N+vtMFZBlDIN+8GITdskts9Naq/0u32dT/
DGZWPxn1LlKbJsgIMazTQbDzLv4fgfiXPAWs60nUpo3M5Rvvvk21JhHLyHhS/oUtkIntWCkOXfcm
YnAmp72xnuNdZqMBHRWvVjbbui5FGXcEdMYIEYVt1hAV/dd0OB+LmZr/j95x5bwilLEl3a/0a9NJ
7U4M1+vckgqH1s5AtGXG+mCLkddVBfFLxS/N+a3C7V1YCu4eoRcAom4NE6m4F7N4WVgxHReAhJuB
rFrTqniz2eFQrO6kAa25xmSUzzJvqdyzhu2oOexPDPr0w1TrF62sJiNJ0KqBO9/Ksarol9MmGlmp
PUtrUKq54tjEDQB/WfTRSx/q4F+K4OB8GrGICKE/QeRn/6RszmC6U6U/5JpeMVD3ah2xrnE2tgXg
E8MT54W2Js2wSqsNo2r2PEHFPbXjFtyKneSt/PeQcbbKSxoFf4XHP6deyu/F7u+jvz4lJJvbnznI
bXfG6upNguhKEfRyJkNaeOnYkGZnr0lkrmxM91tVujF27hVLEqRjTd1ffJFfWCnq5daOt0JTjZbl
tccZXQ6RgqkaQj5ZsyggNRi6P87SQ9vUAcxFSSwMOYX9Gp70fFL7ynychvxLzhtqiI7TklN+Wo7k
KWGNGzZjraYYxsdR6ik47p4CAYTQ0GlUFV6+aSLL1y45InG+k70mqVqtG3vH8rI1aDcVqE5xswfs
k1/yQfy0sHVyohR21ebdb/NJkXUiVh3cpo1Y2ddAbVGhWjHYps6/DEsQ+7h8wZdqQ1v5ugDXCxNU
Z705UY6/GmO0u4R7SJoxzJhsamYXR7LBI9qSpOZtIpmiPohkY+8SumjOzU0KeCUMphPnddLZ7JmY
YuoiqLePlnYfVP+SMbTTehye7OSucVjRw6HIuIp87O9Yy5/dUgqXjMJeXVhHiQnHo5/xYBLqECP4
uX/PNvRK2hjE02n6dKdP8GyzGAXIdT8IvWqzpD7B8NKm2Tx1OiRyP4sh0VnNRJlrTyvkwXEshVjO
UdZQIliaT2h0Dhk8J31hxpeRWR4yGsfH+r1eTCdwwB2wNXbqJ8Gm/B58juiLsFE5Zj/yOZgp6qoR
2IU1petS5cm8ihska4ABzvluhnp6tKNkoTn93fIJWLCnlX0URBSB+RQS6mSnzMe2YSiZB2uxqMMd
xDZ1zh+u9LQQ7sGAbyVTlCC8jiZm4tLD2fDx954oA8JHRr3Kf3F0ipGG8RxVU2GdMlNfvnYz24H8
XkpirQa5kfNGApYKfii7aT+JlQV0ryGG/td9tDrfjp8Tkjl2Qr1YY3kh5wRlkZ/5JRMn0NCR3FBG
LHRywnxUFcfFyBU1WVMTV6AVCMrYETYdDWUGCdoo6tmEVys/2YGAkt8aaQQA9BGNWkQAKNPFYNVH
WGtffXegpIMdLlYxh6z0Dxa6na3gxbPkNXzM7fO6yzblpb0IIzXLk43DvF1bpUNsiRMAD1Av7cUV
6pilFgwNvzBp9S0kne5m/QmmRxrjSjvc4B79EL6M7zoly+BijR3Mz0os5BadCu895qABsFl1pyLj
fdAHJddCH9mqirBJ5xpJe2PJUnQY3EBTU43hPygwLEsRhldt2jmCYwrsbes/AWpFrBpgcGLX8Pfj
jDhiEW8ZTZHiN1V8W6yyi226L48SZZJmvMqOMvxiI/A/bbBDSsRuyci0nMgOd4f0rC8Vl0704aN/
mtG7ThxFRN4kFuj9IB32FkaNwlFf7uk21mdRkv+xhTMjGS7eKsVwsJqvTUzGCLub0++DWKGU+FXa
f9l8UDQAQiDjrti2Qlu+rKQuSoxncxXcbrWrrnSK3rphA+djI49G+QL4LpCTisPYsY5R7TRRd8TL
h6wX5X68EEcb4PTdTIMyty3h397WSyUkCWTjE9zxVrDtEFetJY4IvfqddrTEXw5hmkd0zDyySr7b
hpIqfvcGaJ2IxHMF+2S8ya378L3EZxKhNsUWiloOtRWrGkbaxsLGB2DmveIRWtFbJpVZHARdnoVo
ccdaBiqNd7+d9x6O6Y+2TnskgnvVB0Iy0e+oCO04HofJD25D4uR9IPoGNVYvK38NZO63LpCNB7mC
nMLnkiAM5djVXTKUy7xOWgjBISLLdgwZvoKJhJMStfZ7+gyCowAOqegcanCIcEpXWgdNsrAivufP
62tBlUCJY0+gPAK3vy5PKo52VWZXWriDVt1m9LcFKQMiEPxGn6DLKWblC01EvvzvmmwDLVdA1jvR
/9BG3hItNB3Ek70n4V3lVblp9/MzuB1wDVYkQHC4FRs7vvwai/OxGkaW9XC73OYEtqYuE8Ptn0Gg
3uezvjvgjMG8AeXzb0RJiNwQKouYks71L2sEHcAzT9kiUFy5C5fflRRvmNEfwJO5IRHfKe9lnYRM
CWPLrudlurIfjN8ePOivSVj9vDHTTycpyjrln5ugvUdoeNMkzKY1PkIfn2i7OrhcoEmNkGoV90FR
a1E38GIdzis4lGC/4YyGb5KkEOaYUlMZMmiNNqJU3bY2WA5lPwb/C4sXMiF/JUUQLIQ9xbUCwrm2
+uPToBA9U4+iF12CdRunDfS35aLwg0e9JCB9UssRwOmSTjlSh+PcemvMeo4z6r7NwGmk//0qQiBv
NxDJfpOkc58CdzJYlyhvrXZCzqdcXMhnDqcJG1NVLtvTOYbVd8VQjk0c7JibSTijW1QtdVK0nOX/
5C7FzqsdYZet1Aig8O6rQ4h/ZyovygdEvfy4ptpfX4jPkBUUaoiQB6xl2RL/4J9ZHscpA9/NC2Ho
7AXKWrLa72x4gmzcxV4j8hrjwpv4gyyvoemb8TFEVpdVm0n4/KiybB1ydnmf+vLUBqcMrVzlzUdn
g7OjJmAuHtGaoLT+WjY8fu5FIglPPaXgCvYA9R2rLwSt7WWgZPJ9OwE/aD+TGkGMsfdhJfLiUrw5
2/nIi68/eevPzCfz2LckN1kNBybPuFEpukMhdZFivukIPrSuGQXCX8AybFDLotBYaXv0LLLgKRAA
GPa91SOnpn8MmfGADvZg6qSi0tfAmdtCBOb4i6TXRmWmyPvAv0rNXdInnCR9+c96ZNIdVOY8T0gL
CvpImLjTDUE5NFiG2sYwf+TkFoewVXLUqDrXiGHUswwtN1NEEqbABosf8aFf5De5B1yPiSEYikCq
Gd7Ni6AMxG+FPBuWRBM0VTGTAJp6doCkScrZwAm/qdgMdQovk0nYkje4gSeRo0anA2IrpQD/lNZs
UzEoe0s7DYjOdSvPE+n5aAWkpqdp3SzxanABxkm6Lftfhx5dVKsOGvyOUtMyUdUaxY2nnXigacrE
SLNxgD5A5PNYJzauM/BCH+tnenyq6VMgsgsWTf6/8KLZTiVUzKiH02t74Bs8yJQrAl53csPIqOCs
OwByvH485zmVqNXKrkOEUUW3fd262n6ur5Mt7MzabxfVnhXzDlei5Xb+wIzw2G0xlQBLL7kQH6n2
X0K+yWvb7gp5RsWky/0TNli2vQwf/5jBrhG/wtqYB9+297foU86hMjn+NfqUwMIpzp8uWP13I1gb
61cbmkql6RJ319veJl+IOYoT2OpS2ubc25iuUDuTBnmURhKL7XY6sxzlbd9+8JnZC9j8LwTqd7LW
tx1giincFmKvJk0ZRJ9CYetYzku4kFhzCP+WCjnIYkQ3+TpmxoBfrqmoBUSr5Zcyo5iDmMxPssre
DRICnrfMf2EQ52URA8sGhFZiBk+c0rw4r28lwp/vzqtpuMA7u55jInHGy7KCVu3wH504GOQdEm9g
GIGwZob8fuqn1xBIL/J6BrvwxaxhZ5HHCJOykaLiSIi5M6+ZKmYVIX++Wdlo5VkgNWlfZQmZtiio
jzIw0ZKq55xkJKOvUypXcYrYygMUFqqj+MHaKb765Zz8i4pBqcIV614mEbCDrGCG7JktDa5aYyMc
hyNIOzLmnyFJZYPWRy5YLPzcNc2uz3vObgQlAYY1HjqcTTV8oyQcOlXyz/C9GuWu5KYIG0EvxO8P
07/gS30VaF+OtfH6aICAynsk9XNrs1JSj+7RAaqYYdvL2QsROK3xOJfsu8nQJqlJsfEcsOwZPgft
XG19ejQIJOh6sKv8LvOqi075Qm91QJ0mzlJXuS17BaRBY7Dux8Lq4XqTFEAsKPv7lUTHxvCoA4aX
/s9uNQ8Tz6/ObmRf83A+u6Ohtq3X0CsC0gXA5tUSRXsgX7XIybNLIaVW798VrySBHuaRyNm9tgbn
yU02GTGyLJaZEY5vqTGj/ihBWa9+7wXmK5OEGpT2SEDV7esjiHruKDVnAJCQ3Dv27J8iqeVzFPmV
ddLLKG9Fucm9d6kBBCn8ecOA2+U8eZ6XWNCUsu497h97idWUQz/Zq1OX8Ww/6FdCJOQETjz7M7V1
yja++qRYfSDeamGhvnquM/iFLzOLzt6+84O7NU8270u+JjxqlePkQTaxP4rK61O9EIOZxXIPKxm3
PAYUZiwKigXI/PogjQIly1WMB+x9z+891TPNTVBR07jY+zw85RuyOXdErwqE36Yg52GWjtKLOBRh
YwgN7IH2MUhf83I+tZA987/rL3VFrmlpLBi1XzVWKQJwhWRogFPVfRgUNo3u+3tZWsu/Esq6edxQ
u6b5Bf/JOWkbB7P9EmMaE0OJ349JRGri2MxcJbK0KizrXoqjQbHYa7pgq1FsSAe2Tl39zlw3U7ia
0v1NCe4fy6KAvGjFpGCeiS0LoR+tCLaXHkKNkZXUm3QG8Q7QyqUyfcELg8GLiYIRbWwzs0W1h2qo
Kjz3I+4Uth0uRkfV7mhG3y9YOunx58ruG7BSZVFsj0NHEaZ/vwzE635viRJWg9KgXlyD1Z8JSScc
7NbC1clB5Gw4aIDoSvtvCLy91r1k8XnMkOeKZr+NgzYIXVTtyk1vcEvxyipTxCEoJnUztoF9A/zW
rxvoP+tDIR9cScaKm0kEpgZmkDLOE14WXvS7ZyShKTL+wE+CnJPvz8i46Pk7o9GViGJn+qP4BxBc
YuxUVNMqZ9ODxV2L8e6SgG1NAoB6gNd2k02nw6iCk5FVxAH/Ld5w75A3dml9vSn+rGU5652meFDS
TCmEjUifH/zI6COspgOvzQ5L1jM8wcS4kqUn/TON+EgBOrhYrSgilCDPOiFCI/YhkK1w6M+Xn/u2
OUcm+MTRi95kVs/I+GRqfLCyhw92PySMwW1J/1Kh1tJDoJ3bg7/xPO30zBGaMJsDVdE+jnSVdNU9
FnVcntv9WrPKVTWRSqpvKfcLwuoji5rwmSaEk9s5zSDUWKXhdVb2QwXQ+Ua0U2/4K8RWUHfc1SQR
N2TeT+6nAWv9KhMJPFRpN7N2kGnLa6XaUNPRluBvWU3lb8JF6HRhM9SnoDL5ySCtBIjDGHaHjl6d
YkrNpQqYhSELixToQyKmEDtpTSRu8SfUMWmvqiDYmfk/wcg2TrIqDslF+X8aMVL3utzVaJ2I+cqr
9LFXdxSi4kZjxGUwbQQvsWTXjr+bdG4mwk8wAMwiCyFDXlkxrSfhaoNxp9yewQyyag5wjeA41e4I
2DMyzG5VlVxGxmxtDcc4H/oJiSdCNT2KSxg/zbklikRgshD9Sgfzg9Sj7pe953K5+wsme9dcWoOV
8J0dqyxLQoqhleGPcbxIiqgYCPavFfDskvIvlx/npOnpbEcTI1BkVvYTScGoiZUcR2ssjEWDz/ww
lJGWov2ZrFwLL3qXgBJKXaOe0jwCfT36IkxrACLRg+Zc3Tedikk1qMS2+zKSLqE2OcyyWIHGX8fW
9o7IB0rMAV5N+eAM9adq8Wj06I+06TBvppZMQMbiUG23WKIxWpxL7ShAwwSDJ2Ta7p9h/156eWA1
pzt0kAgr/rq0MNjlehr8klgXUdB2DE2JIkL/wlI2MUq1XZW5hyvVJaXAPeXwWGiX8TRaw9jMnDkd
dlGRJGnIceynQ4LEj0IDqio8fkdRso3JZ38kVGcl3qWyZ252t+8M8mSq0KbaNyUXGRf6jOGi463x
6gE8gylxz6ooDmsS6wlagy9xaMgiSa2lU1GeTzrODbAN7f6P+uKsfS/BuTviFZRtw4u5KGCHKg5U
7GCZGfBSffe9hfN85jtfu9arCrvQwRtdpZUon7/A1PF2vYg/P8vjKhlXmay0YEtIuEvQesBo2FN4
jVO/YuYwBRYIkGwNjEfsWCHZKZz1RvD9TWgrh2lGSmCue0YtZjMjT1Mvmu/ALTXOvp4KJxhVXPBm
PNXs+KwCLim3GrjxCu6UTrMUOL7DWa+D9NSj06zjUvnXOJThMJr+N4LaXUiCbWunqksG1lm5gaGC
Ei6lH5mSE98FfF1QhEVwgVZm0E1xVuvypkINDG0L/P8QCK41mdxRZ9nc6HNRXqF9xTibdGasoHEW
Y8cC6rdG9kZFElwVovNelSDwIamxNnjbaAJ7CRle5NOZFeK9PwX8VgLKUrrzrvlm7F//RpEc52Hy
kWgMxeR5Wk9pfmGE0J3tnANGKGY3igmVAlhsK2lPPivflSoMM3JnoJDJ4xmsFSNVpj5gpOZ//eSm
Pj+vucl4TTr7QKeCPWs89IrwOR1Lt8CTcgp1kadk3jeoLxrfP69KthDGL1nUIseBgJTnPe5L/LxB
VDqazuYAeQYL2NSpYQzmHe+tBpojhhVZWhBp6/AtVym5nftINfhzQPbYz4tlV5P4p6jD2IQbjmGB
gLUhPgE/eCLCaJ5tk3Z9gcR3Kr/k7Rn3yb6OYeD5tbVA55SKq2zxx3OejXYyd7HhYVd1p89a0yod
zK+jjnt26StjrwIzm064MBxSc3xTBvFO53JDXgRII1SJEGlQYGJZ1gIJHuro18Z0gQiPSZznftIt
PbhqKTq8bXHGNo8hfagOEFo1qECNzt+FoZ57SD4v+OXPJsgSkyqXQyMaPCrv6ddVhl/GrSL9oATn
YvRvsae7wpOPuLjKrjmlyI18kRRSDM/ng8bTuGsb7z7nOmUuvHE2CCcYf5BF9U3EYvUR+KvRIKid
UxMJ8Cjd+465AJGtZwvppmLx8K1qtJfp6U73HwlOT+VsOuyLCRvHdopJp834nk8MQ2PKWLSfDUEV
ZJux/iBQeB40kJ3oXrtRFsg+5ncApj55z3WnQwsNy7XyfJc1v4DZg3YrT+G/XGvu4KizmnirWv7g
ydlIaRIoqjPhX3uDyzhLIDEGY88cdXS++PHSPiJsc6O4wzZ485qGwawsttZtc32/5nqM340Yew2/
Ph4ZYyc6wuBsfkwBVsnmZq7MUfkCOFoj44hahq8SUgJXVKJZXK0TarC36fHjzpnyXlDu4K7gZGwA
rupoSpHn7jmKPxQ/kvvLtv3OQix5uyiAnFNUj/0zdKdSbpmCTBPzkKspPg/jw9ItO/lM6Zphr5bD
yZlJXPtncnMxKm2R1tqzp737HJdHPO4hqFnc9eXrH0ekzmCRiJFEsCvcQsHbFO5QY1Wj3oWO8J3+
TTbqaLlF4NRHlN2Qf7KkK1LpGNWYvzFEYUi/kL49UMD3szqy0sPxPUpargRtCXnhSIuez1Tmh4tS
l4BHovZsiWWHD4h6zTSprZO1a/hMoIyBKzYOsZ2wm1U7vjCwVt0RWyF5E2pzP22lwPSrwgk2/PM/
M1Hm4Pl85/404oyrKS+kTXy001epN+vpVrtUQzpYKDPEk/kNYQU9PElMLxuZlzP1CMh/vpgFt55f
bB2YJZYaoucSQ/xLKTBvCm9sZ1bT3D0gps1d1di+SPrHhVEycvI2y7X3R4nHadz4gNkhKIntbbHj
gIHwxlTcFcW38yXW48W5rXv+XQ0UBlHjATUaM5nPEDdSRahBhWPl09GyoGKW+LHc92aOiUhyT5oh
K2tAAcQTnKq5WI/dKrxyqK3SuNwK8AiZImsNmi7b6Fnxf0KG+wuP56pe77mWeQVplZZn+ZMKZrPQ
wPNxmee82TuXqayq4PNRDcLlPSoZ736UDNBZLzXjLEUXsYsOY8BOUWRBZ1asPXY/dTgtkHR4rtrg
PVJYTMPXvY69nBV5oGENwhnYsJnJcBN1D4zu9zEOROJla9eOb3oI/zihgqSmC2rbDdqmD7NLhvsR
rtikKcJz86oQO1lW/kbtaaXaeD3GJg5097oQN4frPgKx8sFCYHa0dOq0hEpHi79/+wPSnQFs7zIS
TMgB9flioYSXCuam5zxKabFWJYqMdSza+OAEYlLBcbi0hIHSnfuHKt4JFX1i+OLKyF/fZ/afc10a
ObWLgrDpbUWE7I95Gng4ZCIQo4rUBve/pa4jrEdI8CClpAtMzjb+E5dv1qLxMxSrC31RpT04lUFS
IRW4ElS8WxZ05qbYVWGen9ZCfm/fVd8GGvho/MFORf4dSdSG6IWIM6QdXr6CCCr/QHzfEnT7kBGF
/C5Fzka8dQ7mxgb0/8ASHGJMSFS17Mpm1CgXkzVAembQqJu0wIRFBhms8ucGRT0nSBp0TBpjvnyk
Unvg3QorJybE9Fk93WlOho6co67vrKJVSwL6rt701PLJQL3ujgMTiJstRoxFH9PieleNsz3qUj+F
laQOkTOgqMY21fB6YHFCqLynbiyvHqU28vzm4wr7cG3L2e7N2wmMermU7zOXMslCKnVu/kTAsla8
GywpS0B3b0gfjSXh1m+fiMyHUPWxYcTOEHm6Tyv4XY1XPZzYLuWQTWuBhRpAINhRq4bD5xsKYBSK
fqbAw6wJZWDb1EEL1nKDP/ko0Rwi16drDoYT/ltIIx3LuXIilpT+2Dt5DPKSc676IEYnVC9sNcgV
EDkef9/j//2BNq+zFBNIlPts56UM47mWLspBdS7cOiYUsv85mAxGrf9grn7z0pt6iECzjmPjIH3/
Q6Yc217bnlczmg7SdzS0Dd1bS/qsOh8ZVNWUU+vJIyCqitiB6mMkCoGF4UJZsLU3IsP8D/NygdVW
LY8oRWB9d+6e4UV2f0S1/nJN9a7Mu1lLDVY3ei5RUb71reyM3ssT2aMY7DWTTU6zxGdlgG86+U8g
+vUG8XEFexwChYA8wDUNVgGQQZXaPmHQhWs4Aw6GYvlGRVpWBmA+uVhMPS28A6uznFLJ+fdu9366
tFjnQeP2vOd6G5SKDNIGtvXyDvLcxGUWfZ6JwNxXQ06m5rrZPRjnRWNibI48p0Ur8SohdClYhoe1
HIN57CzzB9jsTSsy8VfQSzx9Z8F4S/cTs8OKSg3ZwRkNMvHxYTMOMkb5WTMRxhsi+/G585N5KFuY
w+AN9Pve0qyGGmzDv1AMdpkn6rAV0haMi+u6XyByWBoV2zVRUfuAByXCwSHjYSXFRV1VzJlmvihC
N6YqRHLacH7IjbKzOU89IjQ8Y9xyetrZzyaAjyX9vsB0VLq+J2a5tm8eI3SK5AxBp6VGCcqRMWtH
eblX3Oz2RpgifaJHrmuTHZkfozPIXss5dyJOtQNr1QytH5MpGLjbC6fsOvA9HUAR93GeoWcgbUXH
6Ls0KO4LF52Euq0XbjGcR2omIrPj9fophs/Lm1oUypo0i6Mu54Ib73sIh7mXhhlz3ybo3qg4fcpH
ApQEihbTHADhuFoA98EOIkAhUJ1mCx2pQTwM/rx9w9DW7ofsaXv84PTyJMnKXFzvZtCKRJjW9frO
PakpOpSdbA3CoHum1MYr9cyZNujyPbBnLHmqXah+ItSNwsCOMXmIJs98c+TfHVYKtE8xEW6GfE70
m38KJ2r0y3oNiRfUmmlM9EpYl1MQgIsvnb6THcS/LZxLNTtH/U51MNEBxcE54cfbQ9kt/wJiSgq9
tOEONr7oLzWOjia7e3paAVnHBXg9jg6XIiojsqH7uUOrom/0H0sNUUkb2kCvTJBUKOsSpGrTSQA6
aqFL6bxslLXq4aRyKYKcke3Eu+432/TufXohHOZ4BODtbeExsn/qFM5aLbigLLUCjvm4vAU6BsKT
W04YJCEgxonSC25k3buWgzyYGdIx0tlkfV8MO2rKRW1kiDDu0Fm0YS6nnDho3tIJBgL28OHF6dwG
zOGO/sf0Csocrej60dJsmFg5uW1hTqstZmoX0Wh5mZ3qw63YjRzU4gFymkGOYK1ek/Sc0lHawxOz
6pxQ4BedtlhrosN5Zz2l1pGYecSlIJMfbZu4fMwjfQKHbNtJN6YNsC2GCWl4wvLNeqb0FXfxeQGK
Z8x9IqGQwDL6LOMXaN1wFn4PxTZGuhEDIyAWT01/UCKWAQaQbGG5mtscBr0WOgpywbKhh+/2Of0t
qkSf8S1oaYilGswJRGCoyOgGKlCBipvoNCuuWVqB7S8G65v8nMzIXbE/Tq7jDR9FUAdsY7b5rOsM
l9zi8Y61opknEQz4k8ld0v1Bi1igNmm0W+KvOZNl9WnKTc4QAx1tRVAzzleq2lh0HvSBDN0iK4vI
boe6bbz3N9ObbH6hFbGYQDQ5kYX83FchfPDhLU3cEb44DNduSsbWMty/Rg0oEZQ0128ra3BqlRC5
dGKw8KVKNGTMBRZfIstY9ND7RhDpj6buk1IGvlho95Wz1aPBd1lTvwHESx0jAJS4AHDTUgpLd86E
rvHPCYuSUEtGjfDLn5Ti5S7f++nuEW8HQpFdWPToOTgrDaISCvbKbouXYfnVLFH+3IO7LQS2E4N0
4rf5tAoRePZoODrZhrFmM2Hr0vTm/+kyCyLw7AjK3Gj6rLwt0O6sXy1BWf7asY8LE841VfaNzsqQ
z/aJAEpBu97QQ0bpyArtl73vQUtA4TE9xIrttzqywcaIxjTWX2uSqfMP/4uUbJDdBebiEH/TpTGV
qxzGrPR8mmXXuzOtP3BOCmpY/dF+foDtz78nNYrhmbXhUgGnDUH6ESFzndRKQCtMOB2ZS7nJyGZr
bpBWHZKBSMC62uaH3+XE14MwAMTBB7BsK0cUSwEn1Rqkg8mlJwYPjNjMgxT1TB7yjYi4qgUq+XyF
MTaeS0R3zTQpUnfL2DwhD2QEsD0Y8/TQnIUHX+q5zBFXee646/BFK+y/Y8xiDShhtQNpIX7lHl34
Jc+dohIAHrhqskSBJEQkmyCY/P6HV212tzSZIIWgsmZe8/4zl4fjrtogtyR8fktVLSvGI/PFsxc2
RT3GiHiHnsfB4blnpHh6m028Cx+i4SPZ2wuUNRrtPApnVzZPUC/hx9h5G7mM0j7O/M3XvJCZLllW
fQArOYONiHcv4yopybMnSS+eca8jLwVx1R7WNKo0CDTSzIT5VBcYMuUPvSnLQ8oPKtV4F9OkM26z
QReBSi6x0l4WwdZJtxEnVc7YiuuqAT9Ga25ogrjRoeVjhw3AkC/vCy8IiYb5pGR0tzPWKekfiW5c
lp6wiEoB8zAR5MO/34ZcktwF/3HM9oZIxOgla5oU/pgn9wjgUUTcvrJFWH3KdHbhjiP1z/btthbw
c99i7l3Hab2WBpjMmINLVOwyBba+pBmuZdgFGcYKzrEtsp76Z/8ZyToVlilDNPf2QUpjPJETQ96v
YCm5plXr+xc3l7E/x9mj1UlcUCL0xrFd/jZmyHaAeQGRn/zQdjYUkjD6f2LBBqg7oeSh7uwy6ESF
DTl7LuNqXuBuRqrm8mIcd0wNgojtilX/CaHh56v2RvgiSW9rwDtJxMROCZRmb8KsUeFfODs3YbQP
z6SFvDVdoT4eePk+pmXCkiWnvuICDzw+fy2v+P8T+jPwTXBgdVbf/PHGWhT6HfTTSWHhkvNRHyf5
lNlrBfnKhuzVESZlZvtaTVSSXIdT+shL0iOWFdSYg8KYVd79efofDhOeNLt4JzlMk+mOPBUMGmw7
XC55Zknb7tfCSql4S90IboNVHsObkVLhd+XCnSGQTZ2HBYa43kijtKOGJVx0uXwH7ncNcOPZdr6v
vX94KOaCB64R9aM6HaljL4ppVRpb/fduVhuaNLQk8okqlPbRN7PR6nv0IgWSThixQpLMLR1Oqbwx
XKlCFcxXUc8mfnuVi6Y0O3xjm0jS16bQfIMKUZQXf8Rkr6oFOdLdHb3XmhQXgFUxAF6oyYtTWT+B
A4lKj0jSoGRaOOlzuUj4rVk+3x6ftUinttgZRNBkEKU4gN1hDMmitMO8g8sHE3FSoEInrH35Exkm
w5vuLzto7cCahyG+6GWZoOFsgtlubZU3WoY+J66OIIyrmBIUsjCxBPz0TTs/H9uO0x4APzRc2BCt
0FgSDgP4Hv69OhDihw1TL/ZiN+QaLFg/ShKDtzEWdkM7+C5xD4mCkpX2BRIOU9ef6O/D/R8HOqah
Y/yJHrZlQxLQxLJlAEdoMPVtRoc/HYupYw2qbmey4FHzmBW18lRFhrCIVEYaioKb7RWTokI3mNpg
Zio0UXEAf59i0RFqKNFtmC8TIfUNL6MnM7Hm8d6aVRPAyADSSSaWRTFmY4ofvPwXTnHgQXh3Ga5S
sxMIJAGlgR0O2rCEnIT62TigdMdrj0WSy8A7d7hsq0TipFrJEwiMsOiDUgDkiZzH2sC/qDz1nt8s
npwkSrDSbbLYI8JsVvO1ccP65Cn+fq9u15BBboQSzNPWWrAacOh4YDC0WCFIwrWyB//MlYZXA9zH
p9snyRjSrMn5kYB3/kQBeF9pujG38dAfydjfLR4jOp1lbhPsWN4860jXsvfAGRFYUi89esCI1bHR
KcKRmvtKCqIuZZUKbaPlunBnne5IdVm66wTDlSlr0DXVqnJ5DYT0iHmrPjAOK2R9RaTs19ENzfih
zix8pOe0J/G9gFWAgyOSkEsUUw9Cx2tfy8T06gD/rmlIMTbls6Fu33KBXyugcmATwcMCpgrn+Hnx
ioc8rlOroWkGR60ED0W8TNE9dCObEsG8APr2hDBI/JoUfcyOExVR8BBzy0U0fW97BgoUXhLz4+vz
WUm8QwjvTo623hQQu6Amzs5+UwTR8PvC/cfkHau1+nUzqNv3wbAq7NvAEqtCz6YxeWfZ5EfwTUx0
ZO3RWYbGSJs9yLmJ++O1lsacOtDLNOs6zr7h1xlt9Et8TcrKE8bnru3G2qBiz5PVMuNmo7liq5Ai
ceBRbdFbHBPq/3mG4ZIQpb7OoDgK49fvUYnSR3uzDcxcQVpQ1Pji9tL9lVu9NVW4bWDiZ6NyR3hw
GfNq86obmBz5YXSZvHhEYI1mL4PxsXwXPQHNUC9fWusho6T4q+kb0fBiWjxdOMY2kC/ZPs0T23qJ
ryldVkAaNzZMP17gSCu+o7OZpExotaaWF0Wqt/3XBxdf7YMY03VpBvjl4pXhfdcVsDPaJbPrEiKU
XeoNFckBLqfr4eZA8HyeK2DCt/UfvYk69Zh9VaEVDv7deTu9ozRYqeDbokX7AUEr3v6hZqlXfhpf
N+dDeIbym1ZfUWmfVsxMPvkZ7ZJejh1lrIl8oRiFPCIJCoo++DFF/Gx0NNl/zhR3v2RehBag8FBC
KSNeTDgNBasm3VQw3tr5xSzqOik5byC1N7klRANhLTtJ/jBDGQRI/HeRPKQNf3GO2D1VEY/w+zoV
pM2QlmN11EEdig4/68TT2TxYkKIIydFpOinX+tdsQJB2OgNQ4M6/WUCZ6o6mk6lDD8V/P52MYd6i
onyNyXUNSmiwcPexyukKVM3PboMKzMk/m0U2FaHw+rEydhuPlxT7VFWo+7xofcZBkOLnsSDlgOWS
hWvWUVOSviBr/luMyDuEd7jpZY7w27u9fmP7CGIRj7Icfd7BS4TrZGlf5fMWaQ0B1nLOGLXMYpYW
baaxso+a5gvOE5oVDu42mScsaKJTY+sPgxjh/7J04Mrif/nCJIDkAKRB3/Xqwg0kUeMyPzg10ZDV
3MCACwHEmZTZGk4TCym99W0DlzX7naGVfzwSeIaGEanvSLAYBsAU7VY19NiVf/+FYIdPUI6Yr+F+
zDmI6k4onZ9+OyKgunNMmA8PDuGmEc+qSpZi4jq/U0X23n7XoyGCpj+9eJ+quSKSw7FIE3mU1QpB
lXO0FsEdJENsO9Iod45cviyGN+51KoSPITDiwUGndVA2Y7ClcmEgEuJM8MkmcKSfkob+LBmLpLWr
Fiy/jMzZyel47LJCVe7Z9YmEgUbcPljHUFaaHqVWWKVYe/IWiO0FsdWCobF6gCSllwhI0CI7EGAs
ew24sUv4Ui+Ny0V/RZ8dQalVJLVYVOCfAuHbHvClNEU4XUE4reY7WuWiIL1tpQhXOZM3Ihs4mPMw
bkj39YipXV12s2nMfb7Z6rNrIENTmPfBS0Sztz60CXZDKPJcpgbkU6sdy+jy1a1DENP3Lk59SdYY
w3hrfj4vjCI3TiT7w5cUAFGkOZ9hk7697RCYhcfe3fYfhAXIqjmvvPhNGBOcT2hlwqs0MNLKQSPI
FDNRcGtvDgrOLgs4BBFRnQxAe7YV512md7r/J8tRTKtIHfQwC7TpHGaRH+eYGWr1rrB4STc7rx6a
vCXjkBsCPW90cvOT9Xi70FjOGA+y6gADAkOjpX1tkvYMsBR7y0yRdFLRv4ji9gPLzpvaUlGcBmoD
fhC7N9KotUUWl4lWxy/H8UN2acxbgNjuY3M1trdaN/IAd0pThH4mboTw0Y6nPlb3CYaggAWOJLQa
MaSVc8akFG3pkNRM9TW3GF8GmnHjsu7G7KLKe8P9x5VwtL/X2YySJYryeIVY89DodkphqaK7ixQi
h7rL1oJINu0d/C8+/WLG0A/UTcIlUdcnZ3urrAw4aYiOpxH66roy+CIY3qcqShUBeYQcpYPyx4QX
7jrqS0yFA2LCZg8RhZhZZN9z8W96VfcBwVe3g2kp9WtzxGOMK9BP4hNVZmYF1kLgJrxSRl1O06ME
XAT90rcPtn5xxT5Cvss1RZGu5ihKgxoT2mycenUpXYinkCKKIvFI0Qn5uVRQxAQNh80mt7LA+KYh
q0EeBpsKI8uJzefmIIREfQqZmgBOAzxPF9GmxUpgPDukv+JRhlHWAn7OUyyRhypAnLckNvQQG2UU
m8OsSZjZIZUM/w5chvyfWnJYyj2cvpRgofmuCfp4+KSHXugBOdgYSopGSpmJakBE1+oU1ge+FGXr
Mo7Wcv1M9BvvvT4EVwvz60E6QdcR+xWIQppLx9dGutxfBaSpPifopMVKJf2pq+TJf/w8UGcOyA9q
kMA/xSHE/128eDdIeH0TqUkIld+ciqKhFIwjFZGDW2x0fiYS+qpxBxFW+D1kjfsvp72+tlA7RTY0
FFMRiXIwLad1RtTaI640HZYsVGH9m34WsM9+SWVkAXCQLV1HcnZYCsgoEYRbZLYE4bQnDTbVnGr2
A/oe/0Ty7TVFe+QS2CtJKKVuEB2lbex9sobj+JFvfZHljx4PLaDKsRnE18GfkVGYpmWJbMRSossn
e47eBTlFrriuNZNu+YfC1zDKwzipft7UijrEf5r8tsztCx6ageP7mvY4C8/O7toKCH4LnuiUBnZ0
HscZIf5i24K1g1XY5p8MIuK8yHwA5LUm59miQ4l4CX1TAzpAnsmaEhDZ1qQFYsAB6X1Ltx6+MdJY
1RLlcLJ8G1mDPMdMih1QkzZYPVQpc3uIgWcQKi3OeLCRvSCmMN/2ZuTf83KZti6BDrNzMO3bOcYV
zz2NUzmpMkkbDzFxbJSkZIhkYHFShAdoL6+tJGwvzpBLBl1I5W8eevFLPdYd01swyHe9prLnSzsa
XZQX3m8K2h0re+z1/QPtKuokYa6SqE1wID1j7BxV+TxPwFWcl50lqBkLs1vazCsxHBsJKDNaLAth
+1qyipMfvXSB8X1gkg2gXZAFvEj7AZGuj14jMJ7nXz4nPKgAl/WIRX3fj7lilSUKbW57SS5kb5xe
ePVg5kDjgBWcUGJKJQu6TrvHthFX+yEm67PuQfAxDqWbQPLqVoIINn3iBiWFM/ODwVfVT1aoq5e5
8pAl0kbuavyHw4pJRKnucsVUG2DGnjodZha2X0GGo+UGmmBWXyskYUUUIbQT+I/ISeKxrn7VvpAg
/9aM+inHvUx12/1ftkkLdjMEOlHj4NHMTo7zDQ38H3teG6ZYOtwJSol2n5TEsL9Q6fu3wNni7cA9
8wEbxMsraHwuhKztF/QWLF6T6XXZXHoLTHGelirWjQGsyjVukII3KlNu0VGEQ3DLe4yx5BgRpKls
03o+gve12fbqF68EgdMqr/5zTP+tk2Q8dB/gS5D8fOKcIgM0T82zNSUAg8fpmXZkakDb/09gu2UN
OAYuIYN0yY8g30zpx7Ir/lV8/Z8U2gGoRmxbayy0HjbcZLJc2Po+YZv6oSMcmXQeGHy5vbl/6Ko0
WyN1SKwGVsovjYnUbFHiyXEYKZf517nqcf5Fwr4+3UF+omdOIJGCg1IzyMlzwffRdvEpiNzizOUB
qwWxcsBXVNUc30wkWuP/fSUDwGF5Uu0UIHSuHPLh70SieYgUsSggQv1f9QKxlaRKziMxI+ycmX6Z
EEkKHegO+P9QpuTcFpx2aJX3dJ4Ur1f0SZK7pu2Wo+KZYdaeqUUUnOfGagG2
`protect end_protected
