`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gl9vsdkUGsW0AZmvC2U/nwu2OF7f533x71WkmGnxUSd4Fg3z+IW9aDthABVKLpyUnpskbgkvHf7k
dfBQv38JIg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hR15mZaHM3LRqXOKAx0Wt5fGotqScOKkYlcjOb4531EzxbA4i4GIWC0N7wnw0zYbGkXpO8ocsBIr
7LR7G61xy5kbO8q5DKX1O07Zr2nRBwikD4nrngSRqRaFTrH5Gi7Hg6Ov6TNEkf+cyoWnQOPy5BCi
ZmXfhZYkuIYp+EybVIQ=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
i4/lkXkiw7p0eHzSheLifif0JyoducTlrfa+HfDb7Ek6aA4b/Dx4dnN7Oy35Sltf0jSSWx2sVwkj
vNDtIViBoARwl9Xljjcrav31hhHH1bh+dqeLC/0myI8SjXoVnsDCVI33d0nSIOxjt8h8jf6fH5Mq
ey6A2wfGcJj9td6Wl+I=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S0URRsY2r5jR93kdHswnPn/dCS8DtpphOJkTKLNouVNXQQE6LGSCh/CiV8WI6Hlu8+l99q4xP4hm
X2aD2qL+A6Q6/dy9g+1I59J9PHnRzu4jP7IRUuqRnURVzVHMgP7MpeXEtZ16ILAZ7/9DTQXy4rVt
Hmh1+5uPQ5FyHsTpz5gLxeg73Vhpyss7YPweBXcZxJxQYFTrOZigpURCLJ2r9d5HqgE1tUC34Ru6
AHj1UwbSsKGmAR+2Zux3KiYmLK+jA3mRDQbAgqcgNY8ZQXn2NVe76S15890cQBsX5OeCCxKBx4QE
XwNNbLo0ygRL7SdPBmeIEQKUxxy5Ir8YbU5Apg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oECJVy7KkZ6qixqQ24OOAIUIq8pmxvfEdcG8p9iAFh9GciWeoopLg8VoQ/pSfoK/S91sXFgh+FDi
EXO/y/zdovx26KmS4Di3bTbJxW2w6eY1Rs6pTz+4nqYl8iyfCybJ2KG5wesATrl73E03Pcwpr1/E
J6nacnoOmj0+coFiim2igHaoCNNO1Hzo0FMSl9Ea+iBPeZKrlYaBp4mNLVjYbTXGohAGmUaOEa63
oUxHgpz4MWtLRv9uucxu7aVTtRJhE5bq3gs4xI/Kn0+3FKBdcQcf6wnhLoyPK/WnUGz4jv0zUKhx
m5ma+Um2bK6GfhYkn8QLZbH/LVD9ffkC4mg7cA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nTvC9CA1b0B52pc+EmVQthOZudir9f7GR/yNNSZnXPiVCptPHypHpUYExcVolMvD6l8/jJWk11vv
6VKa6W7GXJiUsJ4aHRkXaBuRQVBAQrnNU1LHgbGUGsrFfXUQsetLyOsha+SjQS9sG0K3wL57vvGx
oozbiUY5/I0b0mq8A91CHg669BdDKTB27KeAmrZooRslmYvNi5E4F5wnh4gF+xH4gw0Z9B9KHTBk
3jP0LEjsuTGWXewMgMZLokPk9UQnPRZUg/TZkwt+zsQdEJMYm4fbV8gkuiEd8clrqwJ2Ma0EZ3a7
i/E8hDJ8zefd+T5THG0dhhatblI4dE1ha3HDjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 121856)
`protect data_block
t7anuYJuzxgciqln7af09o1gAmECO6YzDP1IWayhtbrO65FpwrvOPx/nBOXe+Dj8pnHS5/Gnu15A
XUGlsTvPnThnR1Gf7k6WYpQUuoQwypF9pMugipQEx3/hZG1JpAYcNEaiipY7JWXCoYgKYyc6QZNl
ZR6/FjtOd844IrcOaW/8tyZ9h3h3U1IG0ElMGhR5lS8M7ZZsd7KrJ+rD8I5/k5L5xfdnRYR1lkY2
ccO2MZMj522otIP1jBT2FcXzauvSjz4L2TerO+9GL3873r8F/87+mUoAdH5SrfyLKxfeqz1rocnS
TdhUQ/P8c/asGGRgomwvtgR4vvQ+UtX+6xEi0X6C+MatC7XujW7ROxEE17ftoCcKLrx9z8a/01YS
0iz9HT+xhfs4L6A0X5pnIfcY1sJ+XXoZQl7XREpc/4HaPZuUbJaUm5Owqdx++Rl67UuZdTIdP7mB
xUIqGfj0RmmOAp6aBjoFFc+XpdatfsLYbTSfYu1vW6mNmPGFcaVxLD1/GHOR92oe1ju1/yX24yWk
gYTGbXimk+mZx3667aMX14lcH2S5XkBcRqK6BIvr511htnjvEijhHOHipYpHp7ZZawqFRjMHlOp1
eBfEoOv+backDirxV8kfz11bQCX02lyaQK8EZBCIG66x01yGrzUsE4WDLPjv/xCQmnBxW+e9K2Ho
MkQ9Zqd8zVk/gXP0h1fEoIO/IeuOPvLOFrljdMxWfE88eFlgscOblt6nv/nMwDshshLgJguXZe2S
Eo2uILYsAv+TAOWi1Bzjkx7nT9NsJtB6ZaMFAr/heO2+EKhX6IGE/4fN2map8CGgDfNU1DRIea3u
Ho0v4WXuvryzf92TmlZMGCYOT638B6vHVFg99eSljevwYjXU7spWk0n5fefbvSgYVwbsgyqEx1q9
dO7m4VXPOC/UVXFn1lMd1PQ+Prf0A5OTsCUKP1E2PVTUEZanXoYZE6dqITJZiTPrCF5QQuW/VjoH
cctlqyZEq2XznkoWCeItnYw/cbkFpY70QCUl0SSsFu6WzL9HwwQZwX342s+70q96jbrF9LR86FLp
PIusyWrFuqEzeZYD20wy+hjgrXiAa1tELwXzY9ZVR05k9muvEOvBy65ftGE88v8wyRDNDsqdxcmL
zMZSbUbURhhFBb/SM0U7M9HkwIc0TzTJRCA/nBgQW8C5QgHyXaxUOc9kSByoL4Ftb3avMvuEFCn4
ntRNz/kDJRFNSnyeb0eM15+zbeJpZmgR+dugLSFjYDzpKH10r1nPV3OFHnZ0pAt/XQBmclu/dPDx
l627oesHpWkShd2L5HGXtGCmgGNDJqvQM99YuP48LKzEcVkJZFj3W9KPObhz+bP1xAangIZ5RSRA
g+2c+ZpgVBNbeuwQBvWSDcCKgR9f44ojJpM1a15H0JTkVUjcu75/YEyaJCQ2V3f8Qyegn/wdiPve
pCZQbeG2Z4iKj9MEcar5mf3A/I5/vF4zXIKKtB9cierbkTk7Dn3HI6Np/HYV8QOUQTdvSesuoePI
OaEpwcazSU8bHNAcLoKWk8MAO0ePV98IYISczXrpsW4baCbDp0U/bCCjII3OP3X4NBKnSThEWWJY
O1lBex82GR8Q08eWoa8M7SQyoZn2xuXyXkBCExt1CyKqMXE5KT3vqCprZMc3cRbnIyEPnnSkk917
0qvkJelr/0KC76I8IMNDSW6n5ogThUY9ofDdsDC6KzUWTIRZYHJoWYjk871SH2XfQ2mSOL07ZIi+
mFt9/okKkfucvbiwGiChsVLiwnHbp6Vlo34xxrd1geTFQtOePiMzO6z2FEDuojYGAcDarSVPRH0B
+DdLOUBKEgeyKO3/kr6v7xLaT682WYDRYr1ESmP0gH0fFEqiS6UZrEcKtFBPgMeymd09UqHpCejH
81mnabJkAkUtQw7MOwAEXRd90v8k7m6E6+XUpG5+5s0CzIikff/MTnGYJK131jsVdD9dRH6Pyq1F
6viEvZZ+ZzPibwAHIG6fcpdwrRzIVWKwHnrTY9TmipAyOQY4US5XnYWOMLdnrRqdSRb1XNyWYW6N
9M4D+UnFebGUGEZGOnZHqopO1B6/RJV12ChSMUAlL25brLaEX2EJgOw5MRis9zct73CWeFRBDcuZ
V3zz0j2nCLSCG7YbjxKdfch/WCI6xnMlOVYPC1yIA4NPN5VX60XiGm5166CR+shnh6e4KXjV8iS3
j7PWhm8b6iMijmB9laJfv6eavxwZP8yoqZP8OxCPW52b4Ab4mtBz01Iwt1ZnNLI1gHNtMCoPVRlZ
Tj95J4rX96RhEdJuX9j+vuhdIGo8UuDmnMl3BkDh07BYHAXaGuvZzwpjvt/DiTMUGRNrqCM4idgb
goK8ilt6sXBg6PgYi6mAqtIhs6c8LEMuAzjg10uhIsFHawYSSZZDi9U1naM1KPEpaJ+X/PBdnp2r
k9SAF7dicRcSWxhMjcyhunB5ts6gTdxt4mOiwI+hDZV2lQ8TpDq1zgyLdGKoDGkQMH7QxyDT95UZ
Kpj18BC35priVGzD6TzbtYRf63Rkqx95Z3J4Lb8ApeKxoTwHUk61q+J1p7pb374fjzxuK+g6gBSd
7w3n7jWVryMJaTwQII+cLXv2WTNwHbkYCXHtVkT3BDXeNVLzXDAAzk+19/4Kv/ICXwoPj1bopgJ6
chEcYcZXzVwb9fyRmu5WEF/Ld4duamRRCiitUrRnBTCe7fjwtl1PRuyKhJSMtho/hBNvBES+ysXL
NZD2HrYw3Oe7rqxCIBCVxZhLmzi5ERjETL/AtSVGB5tfDtv0s5x/cTx6IqLgUD13OGLRDKsY84CE
+GEmRZ9D2nC08unVClHv7Nj+xDmy58NG+eVfZ+Hwc86aDv0mPlq5UOWgT4R+JYHggcJ9SSu1VWMx
0x2AsLFgrzXJeWAXqoyHojR3rommYDEWdODzgLKdX2Ml4n0+NGePwpuSXszAqm/9b88hNQeIuvEZ
6h/7zoc1tbkK67aJXlh6G4jEUV7R1Cwu2OUS+Vbgr1ZH2FSxpVfpAra9L4b/X5EGbOUeq4DytNN7
9CJqF65frCicOgq1MCqtYNydRAlF0xBmfgp2D5GVVbrnlhN+1a/zcN3lNveIYFqRy+TE4Az5jDTv
r/E4xmBPcXtQInIAJhnhMsf727BPNM51YbJ7S0qj5PfUwTQP5vJMZVArkeuavXXP5ZcrEf8FbdSd
UWlOOOkuTdvLAYS0rkhGSEwstXmpR02AybiDN37ByI5qzWmJujyU0RrzbiBhkYQaAOtCLc3YoB1L
Ga6TuhVGdIDxRxTo33CKGklj7694K3TWuZmY9Ti8Y13n1ISKsFYfOa1cDNg2VBDvOH1/+O7PB8Sc
bHd/EMO6bjlsE2kT6c0TljAH9Ax3zbz5YExsRxCOg/U3WD71iCYJ8dNKqmeRtfbIahtFR5/Vy5j2
qkSdHzaKELQcybkWQfOxx4HwpQpdilZXWLYnzWBpawGOwdGF36CMxMLM4a7CEcUr6lUI59JNA+gQ
XL+J/TX5iLmyi6S19cMUz7NhRE3loTB0ekKfFyW7Fb/ZMs1nGx+lVBIMaup13dApYED4P+oih1+y
szGI4Kan8NEYihIuj6DAELgaMRKWaJT5cwViEDW4bch4BISnFj/jl0z44PbArAN2qe3FxiWG3x0W
nq9acf4W4lMzDy9N8ixkthVMsGqIlVe2NH3rHoB6y5R3t/t7/MiDAcg89k2EeQBiVWFmHNdbSC29
RGIo4T1UgOjoBHNMAHf8S5FCHU+2NABI/Ah38IouK728gfMt9XMdrg1xe+lZGQso5QLMHLXcdOhC
nJawJRN1K7c8bELlQd13WgfzKrba53GX9eAq0+nTClNb2RpiaXsByevuVmDix/xwb1FpsCEgGyPU
wpLJ2Tpv9y5BZ/ZLn9tJD4A7QUMPmVfZkdOWVSakZ4Xos+OjvHFq1AAIXmLF6jocXNRS1oCefMFE
LhLmam15d8LyCqNY1PFc+PJpumm18OHc/GFQ7PgJeMlWlTO5GhsXpI/LuUIgzOPgMAm5aeUhQKcV
jzvRakQnYnkI2Orsi1XYHZGA6EOpGkiuX7j9ENLKtfPFFEF1cgQvkyonasnSGk1RynzYPLKYDwVT
XOYTZ+2UA4D4bWHAzA4PeHhJs4NQ71GdiJUvIpZvIEaalm0AYkMTaIQQsMTLzq7Gzhp41ozYg/SS
M5T3E2I0nQCLTqebX7ZbJWA85oct2dn/q5VVD5f5k/zwTtsj0gvcvRS7boNAMvBsO9c4wg7UHe+7
9H7gbXzD6qjXTvmVB28RsQIfOUQkW+MBvXDbx98+1+83LQ2JVTySSG8mj5RZtsKeBmnoY0By2DjE
zr4L140e8RQJtB/tMX/PIfhoBMyEVFYnHShV36sKMP18XWiynqrJ45rkQS6Anrq6JHLS6J8uIe7R
V/NmI9/8e1e1KuKvf+kaq8kWYitpAsx6YnX+1pz4pb5y2yGODuYRbKaVdFheqJ57QzH9Z/mEULV7
EePP4RXUN3nvkT3Xz5KO3OOUAvOuH7mSHUND3iBcihuvgyz+khUqDfBT4n+5X2SjHUxdbgyU/POq
7TyuCQ+626jZGvUz7nAtRVGs38yBxK7ouQ14u2FPjMIleM61fBDOLNaitRxBrTSwWNkCDAzcaJWY
gV3Ry9ht+GBykrciBnE1Fh0gW9BSa7xIVGrHKsSOVbFSpen8DKg193NVCq3Hb8r1MR+HOVQVJN2V
rFkAMp+airdwBszSnG4y+rEkI4EeMkemcGLqgUDCYFApi75ZrhmkXZT7rLtlZPzHElbB5XPEngtb
w2bGCEmIHQ2Jmlg5+ftY2qLzxzJjszVWXNwXhmUMHvLgGpFpafzVrngsaTLGS3/dxoC1qcf+NiOx
givB82yhDB+1GElMQJpYtTmld+g/obzvLMV05dJIlgHbkrhde3PjEdTka2q5Quu0B6yxaEkIgfvO
GGkLZK2QnwiUrT+5e84NG2lXzWZIaqlRjpUs0oW2qYIa1HDDYXa3tR3JLNbMGYVwRGxcJcZbZgKi
zuqXrhiqQJGZSyYq901iSPkN+jLn+I8+qyfWubKZ0tSzXsyrnCh5qC4L5lYN/Yr243v70tPu8s22
UwOVHegYhQ0twbsCTX6wc24Zszt247uDWnQAT+LFD0nO163nt9V8JaquOfnH6k78U04jI7URXY8t
krzRse06mq91/7HQtGQouolmp2TMYN2Y4+Un1xMwJ9cPHWnf35puSAAXi7Q8vyru3nUfrUrakAM+
fIXh6QTF1vA4wlmbmdcAz3KWw3ZIAGCclERMIr13aQgWaVnjCeesZ2PgfO4XePc2rt0PGuaRlhrA
hOrVrGx1XM6iF6vs38pUgY/BE0Q2oryNlMJKmbdTt9ppnw1FqFY8xPwN2k+llw0EUbjLL+NtE6BC
GKjddeHqjMQWhTYQHg9C5ZqFEaC+jK/SGqD1oksSKADJ4OW6Ir69ZQNKP/DCmvqZBCnwDVk4zBwx
eL0a1Sj0thNgpvyEc5uwq/KvGqFwFSRk23It0y6LV1YiLxkRFQEoTu7lkNhRNljOiuzPgg+37TBk
tiuYUMu3BJrIFFiPSo8LpySX9H4EG7qq/qh06aEMv/Iw+jVeerNcjn21+lUnDzAYKMI12BzzY25Z
Evq2isVfXQVdQPF57gtdfE3AcyIPI86qMPRyUu2vEV2XSLuLLBNO4GDyKUamYH+QM8hErCn0i9Xa
3mnPY3MCdQChpRQ/uyDcffpS1z2Scpo4OWrfuHUpws/PH3W960LCRIIjHvePc6Rf2r33UKU+TwAD
M2tLMrB1bUF+Z0H87gZKd4ZiP77q1vLGKFQx9eakVWL3Bjsa0TB4xxHtq5hUTngoUWEZLSE1txp2
CFlBoXe/jqSICXeclRFbM3I/2dBxBddUbvwFH6PktiuJZqssTzchvSfbuDdyy0WUJKoxKgWtmqZm
sxtvvemfgHCwWSpdjXBeRDKrinjaxROkgFlYyhn+MpfXKpBkbJLFqrfzrdl253Vc04yRHXY/Eauo
mUD+j43SH7MnsLQAzh64rZMrqMI+sh0jwAsqaM36SdpTsHDPg1yQVmbZD3tiw4eFlj1Mc8QnuFTo
WHlwcuAdZP6fbNtDqAQWqNn+h122xXBCPKzL6K5GijtlviG0TAY214iThN78dSV0EXGmn6i+d0hh
gT6W7aWlP7at7EDQbZn7O1Xk3uwLIp+vDm+rtEM5pMmaQv1XmFOAZ4WxPncZyZ7vpAPHnBX4Kec0
YWqvbWwA+cr5BB/qZNW3Qkr0rPb/vvKy/FPJAtFPmSQ/Kbpa2YPzI37kpqKVyUHOEHwtcE/fDoAz
bBRztKehiLqPxh6a9tihdc9NsLBKzXTZTzm5Bj9l7YS2zq2GiomQv+8dOia4ljo+vFxiuj22SM8+
TZ2zbTXPKaP0Tq6BzS8KjmUCsK2moKb33fDESQanOpwvNO/cWA/+Ul2SvEZwr46wYJ9n8vW+yHOC
vauIxHbKCZvqmSkSjMIGjtiI37nDVHl9VNYMIdwJW2Z1bhRiyppXarlLMuZIcwux++QJbEVlqmqg
RVXzmUy9Vom5881FGuN1YdNx/g9zn9Lv0yJ9Wp8GAYy3ZyLQdPDnFO7h64uIxKlI+Zs9wmzvYknA
HjJuoDdy2o8YseDYiX8QZl5XKewQQBdAN0HrLOOPnIY6LRfzN1TdnqZqBlKqjx4SQFi/963SmJEU
cemFcdsucsYEGEkioi6sFOCKmGLGnhbPDiy+JZ+VzHc2KdqLUukKGUssK7V4AZLtFpLHCOGf7PVg
Fg/ml54d3GBbTc0D5nefirUzkngbjKGwTbBOgCtGqNYegLoJEMBAP13E8itkbXOswDsfzTNyxsU7
04cASPjmmOzVpm+wqIAay1KI3eNRe+7S7KQ6IxCD6+ega6hoV2ttznsyp41HzQvUZqFu9Tc356EG
8BBDNis/YdjQXRj7tjzhfYeKHqmvhAiMZzO3NllyzkgSg2FUaykTFj76BPYg7mwrj7JSoqOhSak0
1ioK6vehrptvwnIevR/emEsOs9iRT8mgN/CM0KSNQ/pcZs6u7NVQzPzQIHioK2gSwPto52Z2cYf2
srxSKTfRQvHciBcAXBCkqrAkbU6/TVHKv+jI9zMTF88LSk6y3cCGG+ERMbc4D4fBo6HHHR4JMP8i
z3WcHMjP1NR8Z83tUIjaNYtf+Sd6k9HzrkWGZRI05CwbZSjHFY+Umz62eqa2Qqj/EyBy8vfo/1//
YkgIKJPc78/GLneMtJflKDcoNCl9XMcGczI0OMWCYRqQiQ1MgPVNx9DVf/8xzm77VEDaOwMrnD4B
QdwpE2ZZOWS6X7qyHkKASA/e33U2gLbVS7tthNHgevqbmBKoYdLRpOtv0H7KpD9+4SnmWwZTT64R
55PrzPV5qASpmp3e8MnkZfwurxUr8YiTcGa6jqd1VJvsYbzqZS1Ptue/hH+3B/jJ7U/x2YcBc+xD
dlyoyqh0llspj3j1v+5pb2rxr54gUnTDCQdoV2x1/eTHieWN+CJ1l7sBYSFLExncjSSO551Md1Ts
V9m9tGC2+d5sHkbhSdVENexgu9Lkgzv6QsexU0349smNzjMEahyAVtNLu6bciHEyP18bVnkENGGn
9SAX4MIcSLNvAkRYvnJzJhVhE7TvbBeFniPSWtegXZDv6KVjTV5pYjemGBNFW7WP4L2mL6OcBx2Q
B9czv3VKijHS5hHcLP/OKzCFkVBq2aaWE73KMpoCe8trks3d83uYAixm8esik22cnHLYtIHuP1jm
j4/OO6T6i/GBMcP/TJ/SOKa8rkB7wQFxfawW2zbctz1N6m8HXzT36Oy92utOgNPK/TI7lyZY23Ce
SQR21loxCh3TGGX4OgyNWmK9MlkWtbKNOwBLiGUGo8JflCbPT8ROMUH5e/KP3y6dof0YnUe0njOw
OunwGv48fy9nMhGJE4aAVQkKgXJ72U8mJJ4I9CwAzL1KSQwGJrIpkAVy9HRDAcG8tu9CKsgrJwof
HQU4X+buVH+ecSR83TT+RXh405JgBHbw0K9qCMt7bTmKOFPOeDvuIYDGggFbPWGOade+T01w2Dtk
qZbbhaMW7I6hiyOAn3JLe8L5msZZV5bSekTheXOEXi0zVOt7x92F/eGsjkYEnPnifa0NSnrjAkvA
875toNz7HfLk7FvqvUr1AVRoyEE9K0iCRsjl6ueDNuc/7vDt4dxZO3mYD92L3zWguAW4NLJoOZo9
qCzLnCkMe8Yt2dz5HrCTWPcEtK9yiwu85Aag7jPsT2JzGG4FweFM9jMqWichhATAq59xdBpVpBV4
htnR6fzalcx48B63GKil6wv/FGX+5dD/nvy4EPcD4C9FYRc82o3ruY3+SktucuFo7+6yVweCBDMS
gdVabPvjoykdLvQONyIoq86OtwniHeX0qKEIyQe7LaCfkMNIFIbKDvEFZGrs26aga9fNx7ng4hFC
2PsZQN9f73ba4JbAjBCGM+1GX4SDOJGRrGmblWIjQp+V/Ch285Ae0ImFTwktc7Vp4YTIdmQiEXP+
weQqOdJjmfgCbC4lESio85En7DGLMmvt1GXESKUlwqnxXbMUJYrOCK+1oerAcleMrvm7j5PKtN93
zgrVx4V4YohOnjn4p6bgR/MNT7N0E89MNlOUNxlxT01lTuSBfNHmg5mhkcjwHjBJu/PENiHGjZ0N
FrlPPJvkEoUW2Gn2yLMkgvObLx/Aun35y+2yci7gnWVONqDCYfQaqaCkJhC/WIcA2j7U8nYNrr5c
LlQmg6sYsltyHkO41xceEM5rvgksbFn94tfNRePdHWcqa3uWkDW4m8Ndy4Eh3MPl6aTAZ5E3zy+P
NTYEZtebtCnDwPUWETQfh3jKpcPd1FwNFm7KgI1VK5IeRa//4Pp0KT0Kle5I6+AxdjAQtZh9Nr7d
4reeZkg72AVWaEF1BjCE1Iz/wN5SD+rd8cSNsTGg7n19/+Nx9HMUcRruRoi25cH4T2mSBknPfEnv
5iRWvSYa7hao12q17Z1GBI92UH5ezoLGnSYXo6sIYNStsbLMbxMI9DfpVBw/dJNT3ek7bm5h1+20
hJqIVtAArBanYqRnIDmLasbGrndQbMoRvFV1GfW8iwzB/0jcLq2EdskWJZy51RhbSqRtvYVvDmI0
/6dy/Q1nPqQD2+BEBejE92h/GnoQud65oqD8DBGxfAQ0rreNsn/q7AjN0+ckyU2WI5pA6W/XlOC9
XsuQgSmyvLGeTDcRIdO8cl2VLjJeBu5DW04Q4Ipa+nUb8oXzdq9KpYxxN9leEUMdQP/8qL+5+XSs
Ej0BIVXfIVJt9UuiHY6X0V37g3Oj96/0Gkv2VHCpB/SknPcFIdZVOBAgrM2Zt7r7FTIB9a83WmK8
1LEzPJjVXyOjSeomuiA882LWjod1ogyCYyU6lJKob0pd+eJMFcnsm5VgvQ7Y4sq4NA9REHUGGno4
fUNaYzDfUN59fAwmW8ijsvDgzeaVPRhYVNCqeu/YgrY+cal8tRm0Suzw2daD7YfiGJXK4un8XJ06
PPXGW38XdPgXNvTxnIfFW17ewFaiGuMxEDak5PM+0uZo6hFLGydRlDdmAc9Pj1H+LcrPekFZEZFD
G1Y/5O7sX2earzT+J7+W3cUHZuevAoCmmSA8wdF5WdRCh2Ag3RTHm3eBZoOHLwbJ+EMB6F91oiTf
dF/s3PprEap7DnzsUYmnOlteFoU7lJmNkDbi4r4f1oYd/5D8/0bibhm9bDe+boHQxwxvjvLHIG9x
EjEyAzUmoqKh+u/1eSCIyHngSe/V7c5TwCOvx0loUpqEIrTYHHsSEjAmtBBh5uyb85giCJT/IvCO
pqqxwqOBMYsTSD+G1dSEOKGIHmA7/U1hF8fppNhyL0h2f25objYBhIPHkbDKyqyDB8ibq7EXs9AT
O5KKhZxVCuaXpMrygUieDdg+X0G15HP0oedivzRogOptbgpMNXJRP3BkXSebIvtAJ0fs7MXmehkW
/QRjA3MsH0WoAPJIIxyViXi/hzd4L9RnywzMj+LfyM2PyIjfEaShnPaW2o71RlGBL3kQHkKhXwdx
L+XU9p/jHKHLyiKgj4IbBELE7AwUCfhkOZbnO7JVSnyQu9NVZpMMbzCO6hcLyqY2Lz3SWdMrtoOp
E0nE7yoPcoF9pYA63fsrY35otSq94K8OZP8qhNq1maOPcNJfiD5P3y7ZBG3CnYXzJoniX2IMDkvy
slOx6v4JrmlZzCZqzgrhErt6aD8lZKUUpFpjqUWdEI2hglY2F1JXxXQXLrzd235zkLhoiv/ITEQw
GXSybtU+4dpf5XXwky7DiKdiRtlKBzgvtc76Kuf6RWo5oji3ZHntFB9ZOQ38QVR5OSHmLUNO86tx
ebMRwij+KwYlV9fAt0V7HXXWVftJRBDlEY1e+fAlJ5ytRR8IcjOxbQ1O/sOqoCRXXvl5qFJW0oIH
Hs5P1cOSkeETNlZ9F3q/4JA5fk0geSjDMEbt3wALBvIsRW/pFxe8HccIuJePLhRST+6VuHaKM1CJ
h7Ql5zWaM8JoUhiHnnzeexVXutIoeGC++xogrno8FV1X40RfsXwIOnePOQ+N3jx38LYDz0gXexEQ
rP+T7j830WTmFXXsPDFuuAIAn9QckK30mJoayNW/4jzu1Fne/BYWSzSHeuk3QUSKw5HC5dd/OYra
VYdn88x6v85eQ98pAFNS+obuzgMB63rgiDlWmHawKqqiRJZRmGSx7hLl8Uu2lFeLU+qwCUSQ73C5
Pantow0v+Li9L7jd4J09rmK2iI5o1Qe9jYbgESFOLzc5NfQqJertVUawoxzq4kO9qKlJW23b/jy0
ft3dGY47vxfBNh4z2NLiI/y8u99YItaITXQUxfw9whcRV3V4tYBeBv62bUZmb4yMTE4dpqUiI4JP
Bp9cbxZF2vdFq/LkxmWLq5kOwNDJAuo6DTs156AO0RQMMdimLXgD/XDFrrobqdG6tuwvtlMpnBdZ
AbSaoWpjDev33yRp0TZ7zX5LzQpkFhX4LeavX5NOrHFeoV/4JopIRuU2GHg8PgHh/9xU4O5TRaUd
DO85cRotiRUBJqyf6TdjY9oSkNsBzW5cfOZ0tKEEY1I+7TCUBWFSG3f1kPsG2ONyjlvGlMnOuCb3
UfEMfSWI7rATqRXzm1OQl6CiTdrHZpi3JQoehZKOLepLEj1YQQaOKZ26n06y2kK96u5UgjqJZb2Z
mDWUywmt3sOSVaR/4NeTD4/bvFH4EkrSMWPIRivrKnRL2GIZwhPvvY34C/3qDq5G6gKNAIGG9UEa
wnx5TuT6tV2v4ry4SxrQ8RJk3QCL1cDUuFwc3Ia7Q8PQ19Q8nh5Q4YbbTzOnpzCcUmWtIybsrp8V
BfuBngVi1RhJx+GKx2GwVxdG48E0SwmChTMPsvALQttPTID4or/IzF/eu1g6M2ABtP1iYvXT8bld
CslJOFyGrOd+CB0AbxCXEiDM5qtctcobgeB4Urn25Qx3UTpX9I/S6G/a1djdVudHgSVEZDMk++6D
BjYg2IikUcjDwKTZgysNQ+TF+e4JEJDMgzmioVkWNONkksPGMBNQqrLMHgzEjrplCulDwyY8MCVl
NEN5DRnd8YzJUrJ+4KQHVXHNGMcOR+UBK//HxxnBTyOAujwSh3cHO8M5Mt1L1TH3XyQjsRQcHsI2
vVHJckNDSjx6WBbTjrY9nrS1N7P9sP7HZhuO6uIHq1BWy8QgNIXJUhVhmUs9Wotbz7hA+AscaN8a
hqQMQJKgw1W3ZFj154avdDW8BmUwr5aJSS/+OjFBDO352k+SI8wbiHKdxod4OEwltiPoD5o48zVQ
LpfBxGg7/eF8FtDTd22mFZRnW6IBS72iUycwWIFQdgGt18HeFyybEm/u0SsVHV32GqTIOPoBjYuJ
/yEgwIMRK0rPA7nNSjClOAzFoUOSjN6ZHsJ+6l1liDgN/pF7sqLDsaHveet5yyaHg20rgaB67YXB
M5fwvBrrTV+WcflZxDvhYWSgNlg/MVdB0sAj1E7qVAxPYkwZN7ahW4ntg6ekzOtA82WacJ+QJH0m
hQv9NiZ3yydzUuPqr9KPQg/zC7vF1VJYWdTQ2ZtIrcoJbWHQCYh41lcL4fTMxFyHj7bAbB35KSjZ
foSwOd9zeIp4bCgJqOwgyu3PKoE2pYd6JatU+9d4v5evmgaFmd4DJHe4CgKDP4ZwgOdyKU3Qk8Lu
ZgAO2g+WNUT5zh0DrTyQi26ZDAcg5tnGNCQkLNivLqsPRy5VJKBLrIISeQCa7HffqDJGPGtDk9Ok
m3C8jO2x95gMt1E2gq8JkH/gX3xxz9Plhdz4+uSn6UL4edUqo5NE7zx9i9a7HD2GVrjpwN/fuDFO
73QIAfdY6CwoG6Negv8pPKf9fQ8X9G+fEK9jJdzUDlBlW10lnMgn4hLyFT+akERVCbNwbVwgLTKr
6Pzw6UMAzw/gAgOVD616OeOGMaKV+q47+q4G8v0oi/ZtyvyOrNZO+EiNBZt3M3XBjCHv7+GdJMZN
hpokc4aLXq7NH24X9aWtmKvzCrc8F45FsOByX4LnF7fngnPCY18/2UBFHtENnJ1bPY19Odyb3q5w
uRw1g2DUKX7I+oFQcUzD6ajWVY0/biErXDdj0uU4PeM5bDAqbJbcXl6F6soGbil/yq1NvN183cGG
FG46WhfSSWaZG1b8UMhERla+yiw9/jLubHxCmZ0ldDs4BfBEjDBG7dhmvi5sFIKipRrmCZKrIqgt
45IRHnL+62UDJCg120yOrYWP/q2Jr5daKYDDL9gzJ7jwNwOiBprn8dO6HRUGQsPAkTZ8VReR0fF/
jTHrWl11OYUbNbakeXIXuq3QxwXrf+IdVktdCOmGAk91CHTUOPsG2bmzAcJbc1qwE/QXds3NS0ob
FLGUkHS8fYJLnxEbWCt6L+y6cRwz+IBWSZxkMRbSDOzvYyYUVG/i68TXVj9dDJzkuaSHMEFHDE6w
lTT02x47EA4ZA/53RotRixLtqBcEDA9ssRNAa09Y2IwIZ1+MKd8L5gvstEyACQAJB3Dwc11XWVBJ
BoCKyPi9yJnnFxu3vwtYhcHGXXYBTVYoos/KG9OFZXCrOa8sEy5GZaQE+QsCI1668/F7l3ROEXTR
YsCCgV8uJQdRU8N0G+QDoOIa6lJDoN/edaZVnjXgZqOt6x0ZCNz/YH5rQ0NFx8S840/tc2FRd69D
zUBvuLn5zRhoJwMxXUV7J0VgPGkRrv6E6DWh1Q5SjV0lvN6LqCP0mwW7tEQz6hfO3DgExKVl/KTc
i3aPOiY79kfthKCUZ/I230VeTKLg5l//GPQSeCwyE22GTuvApdsN3VgS8nNL0NG0CEAO7hlIUQ0y
Vi3luYyDE1sa2Bot64dOmewXa2Oe4NY6GIH8ywAJM7Ovq4vcYcHx5aOgV+NodBiS5FasqIz14p7N
V9N5T+xGieYHs2rJBXd5WE0toSarD+AYshuLKcDLbWNqoj2dEpIsYGPMuuw8iq+WCwY4jlLt9IE1
FfbsEyigkOoakVUfuaQX+CIKy3lZauQwiFjFExpCGx0+WqKFA59DaeDt8nRq/8FFCRSEmY2TUZhq
JfUMWFBghYRwrV0GcjJfahNykNn9nVNW7szO4NjqVXzGm0Fy9bdYmk+ddo0li8Tk9ki10SHSdELa
+nHWgruq8cgwkyoNPSJ3HB7ExNhvhEAFA8zHs0to96OCth9NG03dcYEOkrxd0xBNxeWKA7JSZuxr
vyGinNVeyfCMsTXnQl3bssaWdhxqxtUeTG+Tz5ehDUwyrIRF2BVc/Y31DNT1V7d1eArQeaR0KV/8
FHc9FEd2tsNRrz/LqL3+93fPnkS+JXnprQ7UXnMhzxef/ygXKq1K+tu0Odc2KWDt2lcCkv9TaGbv
ABqxiWIdMk4crNAxQ/3tgUT06mkdesxWG9r3/aR1+opesXdCd6Tn4wYP5EcSe1pQWU+lw3luv0UB
WOPxKGfeRS+vgBSJv6VjInz8rEzUSTUVhidog/WaUsYYhESd0A4lFWRHogGGs+LRiVsWjasUM8cq
xTpIRz+Ohf62xKOAr5uYaLpX68U4rw3VD2nqG5zzIfNLd2XZyyGDKHwZQGTIdWzHj/5t67Mewi3G
jdGGGKEmFnoQn4fgQc4n9LQMXETM7hLiXpjsQsZwj0PbQjG/bWMaN05m0BAzQPd89dMrsY0TAxiq
BZvbph+pjRLF9hC9K9PWubnMaI4wRKeppHH2R8fzXj+UTYerT2Ibew887JN/es2ZcgsqicIllox+
Qwtu+gJWv07J1KkQ1Yj4bZZpuq2wJSDF/V41cpXP/4XOQBh2tOhCWgUhtiWlNNUJAOs6kl0EgodS
uWP9+zL2T5ztC5IVvIBNQmuoyEcpX1erzI+ZS9w4c1shA0YhnTiQnA3h276HCaWfKp9NousmZC2p
pSOjHhD5Q6Vv/m1ODlxYVwXLIVOsukpg2fNOhoWfyVsDVcbTgsAv6UAN72BoYjhMCkb9EKXJa3zX
XaHoNzOpgDmJiNmgPJEhjUqULMfa5gYlO2RRvd37bFP9aMWPewJcKP3wdlKNbkTfY+2FvsveemDA
Kl3WBCoAHBu9TSz79b551xHf4XFGWztvEqPfGLtS4e54dLetIBRgqlu9aVpv16HkAozf7VZU3Xlt
QQje16BsnKOvT2+v+pGCzYqpmIwZqTse/OyX30kWSN8dktt50a4WZ3My6893d2m+AgCIavD05ZAN
HJlJzTF6BiA8tQUtWkp5vfU764C9HaKvOYP7G8GOLGS48IeBynL4fb1mo02GxzWo1zuCQVCqV9Ix
/+BxSIpziELnLe9l2g2OqCAT0sUdKIvRGraODQn1RoKySQoWWay+eYXYGBEchJPH4Cp5lxuxGXCM
wYHigGOIs7LyJKpUhOYzlvOxC5i35RLVCvhx95G3kh8QjRO8P9Pal3ev6qlpW3cbrVPeMCcFZFAo
NGd9ZnMLftBcNMmeWmWkouC+a0TK0ampGqNyE7FIxRh4WITrQfTIjInLA/rHz+B0wLZnk3NPttQB
d/X+j9xr/35NNvCnBNqxR3QuuQQch0rd10H0OT6xaguuvRslmf1FGronTFeSs9mrArVJj7GaqyCh
n2cqkIWqYx3Ox82Gz3OYUArW/20ImqeJS3NYjuRlMg1GYqVnyDEu40X6z5rC2qqcjV1VUV015Ghr
lIS6UeO+SaBmL1UsmK2dvXXR6qWiOnJYOQ67T6H6Q1XhpeNYWvY3wOPc8cSpzMZCaBRy6cJXG9p1
6N/YuzcnNRkyH/biZvqzNAGKUkbTTwg57exBDKVHwfdcXfY++BSnYX4Pr/L7Lxask2JzDfQDANCO
LAZx730X2TU7fK6gjY9f5coKI7icBPnPBjGY5C7BkUZtlNERoM0qKFw+fMn3Ek21sLxmGrYCcXN3
21Vpk6AnyoqdyOgx6a42Y91ww1fv5+XBnVigo1QryzOJf27KbK1Q5tMz76G1tXlIyqJYFFz2opVS
SHN9KJAEB0Yh4AZG+a30XKUjAZJVzMyqcR8oDntg3ed1cKcvQUbauox+WRV2MnBR2rj1UhFWovhY
9jFtwNx77UBqxa6x64etQ75AczQCa8cK1Oa6u7j6gnDFMZwn8As5YiW2XLr3oFqMRUUdTl4QqN/c
kEz/TpDF2RR5CU35LnHNxPNKU6ac0lBPRRaGZnTG0lHd18SvFleyIdqWFGh+l8/GzymuhWTIuEOM
PUR8ymHXTA2CRrGYGRol8jUi5BsnqFm6dIcvjlL9oxkjcmNW4Wvku2d28kxUIIN4vittUkVaokmm
5V/L3+EQtuCb/lm7NetwlYO9sJq+aPCfGiaEVJ5k/90GBgPDyl1oU2iZTc9iKVUiBzaaeB3D4Eb/
seEP8gcODhTjqOUtcI/3lqfGRa3vONuqmImCmZ7Lu45TgHvs/0laoersbSHW04OEZIem4SeHoT+h
fZOtwZz79UfKehZeiKVr+EvHMfYAJhbQrGp+cRcP8l24TMNVoA7Pz4DK/kvpW6T8x8z5MkJSF9b4
n1Ml+Xf6BUcdCX2Aui6yEM+XO2XcvNufHJwoeJw+uEzwwzbqEb4mgCBUwWR+JZshOSSTp8LeS4JT
FCvC/KDJ5ETJidSSsWVfzNlVnH79Q7gZgX39agOfFYdTjgQ5Ekjvw9HhfU1lM80484hMJINetTjp
kpzseW15XZAqVmNgjLxQ2AKkWyf9Q9YaFDH4jwe8T/XpAFi1Ru8oJr+c663au5eT/GdDB6/6lR1+
eb1digpyUVQkykbwxogFyX+xD52LiHK5t4/3UkzgKHkfBBBgJm0AOGKcqd2bm1UfMTgouIOPKOhs
PqQ8NzlJPjC05m3ljiwEp79OKb4QUxk3jr99h+1SRxT0Cso/E5zkJLlKZm74mk+wChY0/2RwKMlk
dzuYza494sgkR6QzDHWfmeoDGZF0mrBihGAIajplDdwDy1iaXFvwdmB5WHdWirGZgiz9EwJH0GsG
oV3UWlrqZ/3yAb9QP2XnkadgrAB1SlWN505YxLedT14DXcl2jQ402Y8uGh8uAPBpvmlcnPFx6sHi
Q0gwvqhfA+2BBdoHh7SdbomluBiry6JmOGSGLgi4NxaNG2/3R9s//g20HU63kX6I4kYqt3k1GMxA
XU12i86cm0XysPC8W2t1GwR3p3f+YdxgF1wFS1TR0h6B0VmnRkMpxUV8MStr+E4gjHxvCrDD6Ydm
Z+6IZigMtE/WRJ5ahPX1BXRtFsLZv+FGbK0y187s2gqn+DPu+lISyKN95lqUltSljeeC0H+9dR2p
LOj3xZnA73URc9NNX5TBgEqHeSKPGHjx0ujkJqEHHm2M3+fQKDsjWhliMf8cgTEpH6qEPx+hqfy2
VzGVJR0ygleNHPEhI0r3L1gudaIU+kU4p8SuVUKlcHqCzsP0iIoOjcoiQndh2crYfpwH+dYUqSfl
K/TjFodCT7Vn1SyYD+lVxT8US/CKTcghH6asCabre12/xfv2SjfOtzX+mNXqHHeODB0fCQIMasP7
4rEGV/O6fG4iI1ZWhp7K+58D9TEYEL4Ji7soZrUQ2leesbGBhg4IPgD6gda8o9dzzEv/2VO/JzHe
NrDipOipOxdmmUjwho/84ttRz3e7J1uqXPkNKd6uNuSgO+HoxZS4e6Fx+AkOVVYu2LVbQ92AlcvQ
ALqohpopSYQOMt2a3pJapAxIqiA1ChbWH/nWex/ZMCa6VhaUlh0fw8N5bRNimN194MfLk3wVuMfz
qtEeDRUQN29W+1y6sdXvMeM8nSFe0haVWWCd9yCqbTOfcpeByD9dSE8faP3t/LffwEpmMLjltsqz
Or9LM1MPHoVvDkYrz3I4dU++Mk7S+oZ6HeYMZJWlu0UVfX4JLOvTDgE6cUkLrpqmYsLDZunkOaPS
/ZyMzxdq/I81Cypkvb4yRF9LAM0Yfc85LeuESXYb7h1hjp88z+sc7V8h3zfDOqNv+22RU2FDrHCV
xwmAjiK1nzrAE5NzIr7P1SuOPOEbtrM8geOO6bEO2IoKAfX4MqLK91RxWdHnzpqne84I/V0L6S85
7nQLQG0oyJDalPvkFXuFYiZL12kq3Hr27G093goTuIsBvBVRdQsiUU9kfqrGj2cjhxmou9HrJ7b5
qwSqZVWEuQpo85MOZOQkbKrpfSBJwPHPqSHvvh2McYnAI+bE9XvFtmRX5HoYM0JRNSiT7Gynw0wq
+jXuspqHqNz3mcmuG/SIniLXuEIBI4yrouSVvk+yR1b9pao+PJxB01+dObXGx6hJjgvY1GcqWWDp
oBtNq46JO33EQ88K8kq820/nWmalFrHZ5K8dXrs30Mfz3EydFz49Afevcm67+gId4+a+DILuK1HI
Hz1Arf/C/JgB35C0UirkNkDjHGFwB8gSnIiS4JYBisBeeRk74Ao6p2lueHqz1jIuLUiRxMwSi5hf
tBlA0Qh8FLT2Hkuka6lnvbvH+wZfpjuBzxfPgR9qGSY85SCKoYJLY2HQz9exqHK2cXjqnKvlHjXU
7aoFVaXiOHsAyvrd2QKXsja96F3+F2NEQJ+1LWj6cBxOYaCc2ehQ9YKuElQj5j/lNgOc1PaGP6Yy
FXLfJ8vi9bt+8+amyGWNILpTuhiClG49ICsZl4MxKE+QuIrMfyzxYauYMdj7XpIUrPJVjgvikXHl
JLKDLCIM9zJkH2x5i2VaIyaHugm9HeYYSYV6W5oy0llmPJuS0l4irdSzpnQx7cfcwTsoCpvYn/HF
eyRtLCFCnvg63buLeEij1ZXjha/UwljbcjnuactpmkUEHj+JLdEn7BHPIA8hsSR2ue1QTvo+RSWj
xuQMZgmfdRBAQDeILrMXAp89ss8tlbLzQxw3VrGTnWYCamp3oHMxgLyz548jLXdaHdOvQn04oe9b
NI/ndl+QMnqOhII4fL8r/GJyT5AkOqbcLO16m1dI2e6gsxzxBbwL3eBMq6VTesJZgCGEHXWZdGja
2TTOUOOtH3KkpxMRyyM89W0zAmuI6k1arf16nQblfw3cPG8YDlHfIAtGQ4yOQtA8r0g83rkhNcow
Qlozo64G00ygOBrYNBF9yUp05ulBaPNFuTh5WDdkIl1Z0AMMEH3NVNVhBTbNvvSQFCjy4Smu/Ip+
BIAFIPeoA3M7IdxiVsWKgB30PMclxKRNlviCX4CvuRdkQXQ7ht14IzeP3zyYLgSNoECwxXx7U7ic
BtSliWRFAfT4g8ZS2LN6FIeLWiN+6GSXwy0nDsD76S6K+QUR5eFlM1i7CExp2X7UED+r+9O0YtYG
JQeTJ+l30XBwGU1k2Ev6awI9q+TwHwTaiBfao0cMxmyQ50teOq836Z/HHvZfqUtBljKcumygaofS
DhG1mepwV28nA4qtCuDn4mp8dVPMGPn6DSK7gbIgDOW4md/+HVcWaSqCYkAk6nmzQE/6ZYGr7dZH
FjPKqUgiCMU52DfM3gMaN6Gxj2CLpHgFOnjCno/LLCQkzluYWnaVwbMihHeD5awoYE9aSdLL08ju
rZKiH0jsXkPMOmnvIZhGjSvIuFpPbV6niyJ26GirE/UQbpkjYsu383uok9C1UitUjR1bLFinmmDF
JzwCxioE3C77qwfv5WmDRGhJ9809DoM1YD3vGn/DYzEG7MkmwIAmFG6KuW/o3PxJBtMMU/MXgpe4
wt1I93ee9dDvtWGhuF4ebmunooAkzY2jthiM+CeKR95wrPWkooHXjJ6uIsjLH6ZAHcEjdNlBS9Px
NjE5QYkmUqEYk5ljDD1F/aY5iZCla2ZWBx+GbxlTg39c+hVgPlnPoJfiowv0FsndSPkbxneTtiQL
HpsTBc2D4C3w+PcaL6Rm7SLYvRW7wFsokyZ2A/itWtEVyg0JrGQCXYPgqk7Khcjs2tsA0+8olCRl
B44QH0YBGdMxBzJDxGBLckby020gdVponjfWZcNuIZthkbnFaCBH4M/3ngFdK8sfsZJ3PR6evBj/
kq/wpa4LRL0xOQt7lOKtcuxdoho4PcvwdhGgrDBGSHKaZb597Fepxa3DJMTc3k7JLj7ppwo2jg0P
Ph/gIMSCmRq0Z9pPUmd5o8svXpux0I2DlscgzeuUkPtI5wPf618mwmRr0si4G3hntUxItoMw7SVk
IyAoFAq+v0k0+4ZWkmENKbm6IT21FNItTmX8FFPJJPOixI8YUyX869YhYFIP43wCwaxGsOEuaKxJ
j59Rbt6ZvqEAk+uYG5rQA9sHUvzTZ01YDteGjItuIlvqub6fu0granL1o+dy5NJOHAz1hSmQ3R6O
Pj7s4aXdjMTm7IM3nGeAVcqb1jjd8kEe81IvWFgjM3C4bjRfCGPUuMAKBFmYHazhZxAMhuI04tM2
M5oCNsVS+I4Y2EqOlJvEixqf5ywhanpPI1BphIGTjMp5tB7YSb8ES+w/nIwOnnHpamEw9S71ADVY
Cb7kLuzg0Ez9S9woOD6UTNpJoO/2oXOFt7YzVMlFxNyfWR+NdiZemm1TYuDIJiYhyQ9txfxeswU5
t0gI1hwYwHyM7kDqwdoMNuwIPpGLZelpr6hxj30JsMsMCPsJRBdpvaTGx+Ij6SH04OtnSylIDieF
XE+RgG4/HUTwAqW/KcIGjWp9Wmd/up51XofWk9OHc+3yTpI8rMesotqF2/vKLwbxUYXt3HD+hzWC
52aOP/6UryXXDqEgHtQRQoD/HeOmK0udmj6k2hq8oSR/ocHUcWmHmwcBb/WF0+9bjgrqJX1x8qO1
xO+1gmmATzy2NoS41DoLehoNsJwhgM+MFYQyx1UcsbsOrTXfNsJ0eF3VLH7CeigxVanrxtyYj0XC
fuEwWxqPXUirhn0QiSiYruL54+Bv6k0yOuCak3x7wz2jmHtTrXYyM8DSKwQIxoE1W9FEUvOZv6nh
fm28tG5r4oiARPoYnd9JVHV8Tv3JfGKp8duQ77CpcyhuJfxugB1YWlDzGQRryw7LaUc72hPudqO5
1UQKivCCxnonCpXQ+MshOro5P8jdFWThxNiw528jfVqVhgJTgtYRN3D2gnhVX0Yoml7fuuh5oC8m
fhS/Q2eP1JDB9ObHBt6yAQpjJBfOm6oAvabUyQmWisGcliP0bfPw0eFIYB2gWkZvzJFMdA86ZKJW
VbT1Bw87ovlQhxypwHvpnsBFkNn0LHMavcBIrD4ldWXTPaMtLpY1Q7Y3so3gME/lxC5KOJcQF7t8
snPSSJNMfEPLQHlkVl+y4KpbullgYoDPkpz7JvRSU6o0AzPzgA2jOKJXTviVhjX4LYa9+GqXN4Oa
rEcjEOvHkvFON4PRcuOwHIuyvQRn3Rh6acU165WGbSS46JLFd+70Ir+XMeb87L46i1+MiXr+HoEt
479d30nMKcl4ENIBI8sBGGJwoInoWzjA48s2TSduZpICL3CEXWtWW8Nr3VdLbCStTDSXIMMZdjiu
WSj3ycNb5CcCi64WAf0fYruM0GkaSHx7KYrPS8RPJ+nsoAb6KhlmjfJoy3xYNHZfcXsoGrXDr3i2
bQlw7Qs0OuoALUticD22mpj916mODCZitD6nutwU7nPpoCuBbW36uDXgpS3Hao5Bx3F8RgGNKg/D
9m5iVQUYBwI4gLEz/Q+6ggSsETArT/rGMHzEhMPnvDzi70STeQaR+CsevIeaDtNdoqS6cFXzWafw
II4B3n0krXNhfskw4DeBT3CQcLcOr9o14rtyDe2i0Mk18hqe+zvn+LHey5JCYIiFh1knirWlnjcz
RtPv1wL60YxiQakIaWyUrvTlbKrB06cvo9CGdSS4rYDxWUndB8HlcA1ygWm4CYgklJ50Z3plzBRu
d33MlDrPN0Wbz2NPA+ywApyUiraGmblxPpwhI4hGC0AsLQrqHaMv9RDGZTG9O3VTfZz/Vox2V2VD
TvdBiOuZ9BAPCV9zfNO/lDfIzVEwlKiu6XGfek0an4ImCeyhdVA/uAO6KuvvCVLli4ZRwJBjFc0J
5UERWiQQzXo8Ni5XOdz0VLdINwgoOoXN1j7tFQc3O15/gjVRrQdJ/yrlR6TpArhoHifsMaluCH++
ekXaNwYG/ezJiWqHPg7Wr0w4biparG4SzzzlNOpNnvdfkQQ0T7jnw5kdZGWAxdaqfCtJb3kFJPoV
Tm6RCW9FDpKgc73xckFYRHvERdJ1eToeSVPGtwx9tjWzDzozRKTBjdfMlHFOH+R9N/YBqY8+bhr0
BIG4ZcRFC5R0YhYGgHW+xkKrpdU+znHYlSLYn3HA8QOJ3r9h6pUsnuxVKBkjnfakOtALo0tv8raH
2ElIjdpbpDZKLxuZ6WQBkWJvUZ+BhjvuN0cNfhgLLgBu6q9aOH2W/ZYKk6xx/Eh5zYS551th/YfS
7SO2FzB6FdOiX9srtftmlnHnK4szpdd2G6rVvNeaR8hHHXfUfTyI4yuuGqd42SInS1CpC0L6lIwK
CDe4Wq5lxX8HKJiNnGHabGhAZfpH6ELsDvGt1vzjbCTnfkq3Dkb4uj3Q9KlgyvfjZuokGopQXwzv
jwbUMkwthB3REUse6Klv8LHyQRtBMwoUX+t39sg2rV3pijKi8bpVDOu5M8AVTrxop5COG3RlgZs8
jR5OiovEv4sq9QyISPKAgXpOk2AFHaXZgS7H/5zLRNzXv3DLfVs7yscZTTCPqG+h7klwfAZ7lEMR
k0UZVYUV4I4Eshivwtli5LDA28fw68PNq1e6t4kpNajoj4hQIS1rjSWijUPL1f8GUrROW1jUjoWl
nIz6gVwFpxljxRf9U5GBQTFQ706R6ZaEOzfcHJCCGA7i03ikDfmqId9bdoJPjoVkM9PaXIaJDxPt
tLYsUWN/5yJrGEAxEM7LoKLdG2CenNrCbIb8QxHMmo19af4NLF7ZSsPo0KFS9P12lXcBJ1s8onld
iaBj43pX8J/M+fAi3Ff1Q+RRlz/kKChALDbScrCNxZCKXmS7RgbHm1z7H0W/lDpjSEUwcNC8+zoh
viP3IT/U4VAZt2FsNNXCyn7BH6JSLO2wWWMol64hG9ZIin7TXrQOyavxnHCeQ5xoHgCr6J2Nwb8R
3USqPGW+4Zf5ZSeXKeVrZ2TAPSGTALG+ytOhmoLy98CUoSpS5IwWhxAsi/hB3nYl5iZGdG/Y21hj
pUXAUlRzG69Q3dYZUk6ubfF+l2ZfmtNjDeuU81XIAPsLhN6fDi2TDsDFWJ4ydwPUpC6P2POl+3+B
iBP4IfF8FuqNaw3oYfFRW66qsxcLvSt86QvyHEnvG1VrrBkxrLLpGHbORRwShFjMtczGZY30HI3f
YX5G3HLcSYPVWxNNg1OhOi8cUnWrxEZJYQ/Dzi7QVpfQQMLqUIZwsBUZ9j35OXpmhGrHemdNdLCd
l0kFlWNmLZQRvh+JEGXU+lXlIUKNhh/c+TWnbKsx7IfHMVkP4oD25L7xZv6q5k4Zv+cxI0A3UPp8
xt2dqfWjcqgzvG8b4Wkpyp/oaUYEDQZ5LmzADSM82PrTOvgEEfS5be/3YnbUGOcEvWUscAw9nS2c
iDglmdikxtpjX7D4tqnBifsv9Zs2JUjJo2iKrLoQ1BrBnZ+ID4chvRHhJR3PUOd26FOgrOChCtVq
Ey3BVnBSuEGJJ2Su9DVRsJBL7fbcweUSSQVA6anmEZrRD+sel1xrk22dQQV4LEr1YXnk2h2bEQQq
4ZkpV3T0xBM+37ewILO0ZwpgztTI9YEThuuVyMppDF/x7JJZv/70tg5R1yR++UYi7oOHJuMKHiuV
Yot3tevch3iU8c8+4qEPqkNDS5CL4Wby86r0fukUg7vhnVDkC9/jraRaKWKMC1UK+tgKvkTbdroO
UBO4JqsKvHgTLvUyX/rGcJjiyLtrZjdXQH1ALExs3yNfTk3VFZqrvz3rWUCKTKFVg/zTrar4+qMe
N0sbHC0YjLDMS/GjdrF8xHVjbTcITySKz8AAIPOBT0ufMBG4U2oDpH+nQ3uYv2cIOKY2fmIH2zos
GPu8UoEy/MGciFy133AuUT+u2eIrm63WBvH6GqkNMz2PZLeU4q7tgQfy6sFNukdYNkSyS/PITnIH
ciI7zRMJjFbo6KzoFeDdq6QWxPIdVB0Xg2z08boq/9mzpy0ZtJ5pWLFkUt3dup4GGBRdTocG1GoD
fMYS2K73X7RaXFEkMJm2Zvf4CLBXJiJ2AsGdnublwc5mk0TgBfnvTM4INDTPjQxBHqlgXeRJairD
OzzPytMBcf2E5mSe8xKAPb/GLSJot5K9cE1AxakqykQovpUVMTsRh3Uh0CMbbgkcGLREcfasK9bB
XWyHvdTAhCzV7/hg3DMSSxovmVRH+NYhSpH6IcpRfpl/UKYYyt6fal8R++HASI5YcusxBkGLtnct
oejfqgJe3ldFLP2l9I0qFGK/rCql6WToKXwYjylaYi31bDhNCYdtn51dviCrlRuTCdVYAQZcrc4b
Pzyplxk0o8YR8IHRC1pkT7JZxLn5p3z6SbK481gBIMm+Hy1nEqKgGNanz0oQPji1/6kPpU5L31mJ
x9kUz5CsoxVFj3I67i2SzqpM60uh8RxIlKHi4DyM3ws2ceL+VzpJXKYNbt26PJNBctyrN/+zk8pb
YTER/Lsor7ibcmgGkX0jZ6vKxjztH1IHfKptQKO/F6c7ydA9fokqpbpnnpg4x1RaFjudo9dQskqU
yRCZ4uMloU7WDpx7JyuuHFGBig79oIQjCft4mw+5H4W3aKNDvPaJw23rpHPfgCrbrAUChi8siKlN
7zjUi/kFZu/+BPvk7NIx/Xhb5XVFGR/92ETuPiS373nVrzlnvqD4yKfGZj8z9ew1pXF46P329MG5
emwo3UB1314jkXcilmbtmG7zNVKgbSNyekexqP8y4eiuJuZeeJXdtCQAk1BI3QkLFKgdutoNazOj
9VmIwF0+TkFw2PCf/eoEHvYLhgBNR2KhhgW0YKXlF1ZZ8gRaahj5TrGvLFJEsI5YzmfdELz8Umc8
+5ndA4sqeReFyqyoVTc5WxHeSYL3ZAQZSQcyQ1o8d1W8iy7s9Qoz8dNTBd6SCqeoXSpSxuKolT47
bcyc3E8NLfibESPt3D9N5zYQ8seoM/R7BRkJ0IdwZgQATLdcrle7+zS9AzKoosYPq04a7MR2bcUU
JTCxo017tfcuYyTCRVoGqYYxOJLNBOYZPWVsJKpiuxMVh4Xdjp3lXLWP8rr0zZRvMgF6bFFSzr82
u0qMDugmFB8NDcF7/NNQLGDlJxik53Gj/jbOcAmHjUnJM7tL01sPTt/Wwhqb5GmQn3g/K9+diXtJ
DC9lKmemiaIDuOwYQTM6/H1+98jiUVHjXgk5oR8bPyMPt3zFT1jBErlja+i2p69jzXGqmNM6Lzu+
gIHd04BNd9RAk1lbJov1KNuGiD7V58VLxA9HL4Jx5Iw8lAGYCn8aUwIAEArsx0Ca4n+z04HDeNT+
O0GYF4H+bTyWZDsxG+1+Ct0mCfTeYKRDYOKp6HPIGFPr2kGO075EYnbW5RTVX66ZoEmBl5zO7Rem
EF4exOj/twR5iNeSoH8a0GuqkKd48Q6y9EnXRxUUM3BwedfcT/UNzuUj013CipUmCwBzzCZWpLw+
YipcbOrGH8GzMhwsz6nUnZEq27T/L6WTUmcwF6+pRy72uqCMGewuOVaQ/RgWYEbbw2ukMuKf3UuS
niG/bDiyeIekTKVy3ZMqsxSNhHV+zKwTR5Wd1mFlJABtvh1G6xZLr/WN60JMbZOw5CaC7PSjvFgT
l3uRHkR5LHINdkAI8U6vM0BmncP5/UIc0ZN5DeaMTrrpbxOfqSV0Q9ALbI7L04FIhaSEbQ5VMet8
1O6b0el1LXNISNH3iquEYKti3e0YotYgQLORoySegwS2CMCuyr2SHtutqrFr2urvSd1b+k0b/Zje
p6+Eu0+647ehu0ghFETdlk63HDR6mLqn2iFKf2jQSkQlFFyWMkOmSKDnuahb5egt4ZyMyzN9gLN6
Rb0h2cdIP30wx9AAGF/lq5ICKgDaUBQY7OFIyJS27Dl3M5ZmVYqa/pk0HQKIpEGOB+3OHu6xvQxb
526arXO8kU/+t6U6hQEH5H/qkBg3VlVQqjaxrymgNuUEXdGD3bMZguSMj+YkgkKIDX/Huw1tE8Md
FM8gAgRaR6PykfpN4bqxdetzar/Toa82fgEw1PHcA/L8a37iS8LETVhpAgbYWT4GOFByM66KbO1q
yMcidI5zZDKry+hzvB3InFdmPwFXGFzkP3UYQgJnt0xylZrtn4Do6QkctOdspw6B+jxNHNgzhrW+
m0xBIy92NUEgiv7qXJkCcqgYyIJMiJbV9PMjjmQBIk1ZtIY/HFqgJeOYroToiss8R+JPpEC6s2lY
4JoaW2Uaw84+p/P10ECwhOnniiIfEYOhnBpvBaVjDAx1hFhxsFYlrdHMarcoUVhQ9LtKpUzw8nTw
OFtcfw8arOjrOxzFXGcu3ZIv1Xg+Y58ebs+JtLXjDom+R7M6vn7WL4XocgFNxwP/3v6JnONOMNQG
mjYIY0V8G5ALQ49Or9/0u1ne8R52G0fCu3gz8/wi8WTgzPAt0Sj9S2HtQJtUBi19Wdx3RVIe1hPm
wjRcXOe3AdEKrmRllb4s88B7LBJwmua0G857mlYTpa9lc20mE1ry5VQP/R3Mxa7CbNtH6CsTXb3E
u59o+96ZPpouLl/B2VWnMOplln7HGvdwc81R/vylookQYxBfCU0U9vEsvr2UpUxTKFR/ekhbZP62
26h8XnWWhXANqtKgNObUl5vDnzgx/zch/vIHuGd2eRybRRNdahg5VI5E7oLNJyglXmqYfSkS2h8D
llYghouc1jGv14SVySkJD+61jHj91EnZgvB/yZuaWFOMr5I8hB9RR4jKlFJm5Wq6+eohvE4ZjPc6
a8aVMrieNPA4rUhXuYY57D+uWDEFrGZaCljQJoe7PpYJHh9cHD/h8s7MGaSu7ZXOhWcRlKSq8+X8
fCib92xDaYf9CKKIc425n/n73Q5DH5MWk4ZFdIRqHP/R+E4bww2Ad2UwSa9aAX3bJFMXvY+5Hzsj
PCYHbYqLowUSaJw+cE5oa9vpJFO7jPwWSgJvTO8LEpW1Hjc48d1Vy86M8Zjm8jd8CFgc5g4azWvR
Ma9Ngl++eyOsPeKhBh7F1jcNaqikiGC48I5rVTXqNMFqH1A7dv/6ahrubqlGKbYe2IWNlf7dzE4+
B+sdvB+WTOOP9kHni+x9TEKm3r880XjmZHDph2SnHK2JPBm/vBns4wvHU8kbRIDEJ8NWE4BCdSYM
QFYa2TzszRn23spqFH84WELFjvJfvzmGTJOp0ILUZdKGI4BVy8ASPk2c7NEx7yJ/dr7bwf2z7eiQ
9zw9BdOKywBCku1VLhXU7BILvCjfIOWh9/+5A+W4aciDARyNr4UqSgtOeOn5u2NbH2GQewXnQ9Zt
jDRcsY4nhG74BCY90I0Iv7WrZmk+6b8qgWV2TgNUCS+UiZSQrDor/mGvuwtYtBzDHb6gft9bRPKA
J7pg/sH7vffeTcVRFrlyciLv5Ac8tJH8n8E+SytVZxW2+jI6tGrc3cI9Z79Kl4BxASL41MMY1l31
OdvXOu2SZ8/mv0rdyP0CrN7ekK/acV/sdxXdLC5gvG2RQBT49bmbPl5UaXA3GTWj7cf+vMnMq/Mr
hn32iGPaoYx0SG2uHtFUhVB5EHdkNHe7dnxVr4x8DH7ORucRwjGerpmSBN8RW8lfpalYbelOOP5k
sCQsRYaIGCG4lY/AWgFOfmL8jr8t5qhYcXf7U+zaLpxpIBvKZbH80V4N2uJhhzR+GY+mIJgd1BCw
IMnXBd4YOw/LO/UxeXGSkQVV5XBPKL3OVhlE0eDN45WQVS7WE/ESJJqKDCi4BEDHnhDfSBNqPw+w
B2L9T7T0QS8+qy9uTPd1jMsS/zhoZprdHJrsSxiVdGMUuOvWoI6bkFvslJ/esvEJXrhrqi5Q3Qbl
Dl3ZM7BN8/RxJBWC2c6/bK2xQKC0hxAXjQD1OE5/1PeEKif+jUN3/Pyck8WJEDk1R+spUNBPNBBy
MCKU7gJE2SKzHxJw5dLHXSU17Kp+vLB21Zi/3gAnBCq+0O6oOOUYXEpbMcI6l/5JECeh9BAHGnXp
g8tipUCasUk0y+wGuIXxnGyGPftmfERSt2DkldTozNVxkc4I7to/5ov8VaD1fSYPU7QVImGbJcuK
TygfS7dOTwKoGNMs8Xwp1XrVqv6uMq94tv/GAYtRkfR7u9u/286ux9FLMHMsMd2Tx4liP+bEA6Av
ZD/UX2/0txG1cLHweDqaMOewITahXoASQVvr4Ivb0r1oCwRCNtab70C2JsrlC8pvpHJFQITfkXZN
CdWduvQOcyFvXxJrRTL0Lbt7Ed3AQDkjHUgzrC7ITghgJwKUbyaPcuAf+ohaPHeil1Wq0O/6lDvy
i7GrP/A1AVVgrrspdYKlKo4gxH1TcgzOLbXe4CKDjk1rZGyIQDYHyKeR+rDpvkJKHo0q9fGMfIPS
P3rj9eGcSHFGl0o4XGyJ/rSr4BcLiAVrrIYdBm5ltBONF3WMmy6Nv8233jXKyMhwmnrR4254zBNi
/x1RFeujKbYaKJaTFkWR+SNscKrobIDIIEv6TUkF8dk9HXU1V+4Uzbdb5eM0tINRg9NYWqbS58bk
+5YOruFnh5vhiLs7ep1npU5vMH/5BS5DIab/WC6bMdaWcQDvepGlfXLVPXun46hCiKG2YJ4T7xQr
FXlPx2H+JWcJPNESMUiTIK8m/GFSnzyer/Z1wPKiDqVsHwTBi8aowbr83WBRhWsa9kViwNo6YUuy
GUMcQmVgk2tT9ONRQxvpuI5ehkAXvZSB5J02Pubiyc9gkN9pGr5SJh3CqFY5uUcV+b/ogXzaLFEq
ADvI5C3NpH6rrja77qfwMEJoJCvQSYEQGzHVra4/IOxqmtesRgoj91v/13HMonrH++KPo3eUPtI2
WbpWjtaBQlBRLerA7D3A2POwsj6rdMt8XhV3q3pZcgT9EqfEXBIpBCPR7NCOIZAQqnDd2oJfJOk3
WGK+59LguvndSW3W0kboZCEHRTGVR2wFbnPjtuGC32denKmj8bduC+jhDDaplOCIfYDZOPlyQwCt
drekc+0eB0pt6NXXigJK2E5kViO/PGwwdAjt7gnKQ3ja01jaQE37Rnl4yzH4PwAWCLZue5+BJzHt
ofF2HmoZgbaN1WWq45Tv6fu/ztnpGJdfeETRtdioNdJlL5ionX0XExN8KoQI+RRuLNASvx09C/Aa
VEjHkQSls5Q9FLSY6zqH1iAvOA0nZUYtKEUjPj5I+9HqxewZf9WGGPNFUbG5dZ9lICcyGdCOrZfc
f0q5REZdkoLmS0do+C/AaBh+smFLq0TJuVtld882m3Zanxyx9Q2DityJ6hFDHATSHpcnypfDO09a
bETvcdgAFoHWtMX/HtPe/MT51DxYbx119JtcN8WCyVKYwufXfiBGA5sX8pIdCZxqEncu8IGDX9cu
qJN/UfzicmiqOAc4dO0WJ3h04/deGrmcyJrQkm2nI4Xsm2EPNjKDxdu5fA9CMrhed4ZxniJSD3lz
z2J9IcFoiYBnNB/hS8rPrl4EZZgeA5wXFNhlOrPgQNLPXCUTn9hqbMAjN4iW987WKVQ9jV0pcsbk
1CNP/UuSF9uIR4USRimTTy0ZmJXcsJOOWFGKd5QmdVi7nghks/OIngbUtHBUwK3xzp73o3wHpJEC
Ky/aW4lYPloT5/E0knNpiwoyW4rYO8tkpLg1pugp5pajxRG5XiPtSfZSkOZpub1NAqTEN56ZJWuz
iPKGKTktZ56I5e9ImERckzgodQLBMJyHu9rNtbAhcf8WvuHPYNcfVWxEaRK/QAksjUCnDXNXtvYA
Os4lOsu8YncnTxvRtVe2W1cQdGysyeQ5IVeJmAsayn5I94V9nIn/Y4kbh+WOs4SArLYxUSf3I7ys
7502sfBM9XWrqTeZAUtWhJ37cVwHS749ZzXE0uDRQ6fx0aoILmoVOlQx3agyZDB6f3yswNAim3/u
NcSgeu4czCZXWpDYarSY8GjzxjDqiJUa391iKEf7uxGaCvS4k6kZxEyEiedUvipdhOdzB6oJf7Nx
0TGUKNToKNzfvxp6ZOz9eQisZbC1SLAYEN+VISnmi9Rdgq/EyqYwW2Ku7kQQ+EJStFoBfbgUE2TX
IYWo9r/F20BmuJkDqP/EVlMmuPCPtY17Ia17J8pIcCi+caoqnjKPYH0RPRIBJ+jVDjiKPQvsqRhn
dxELhV/LrsFT7R6gaT8B3PyWEi8YYt6iQD9PvBFR1FvrhJ9wU4sn4BZYLCjON2NKVtITy45LoWyo
rXonob8bWDd/R5W+JS8DDwCx5McoyheD954qkqMAeM2hQueMOvyi0bVy/LP7HK0uzEWV/GBxYCM9
CpxxrH+8FEVfe+gaJi0C7iWOCikwXFH3l+fxUks7tOi1FVLDlSKOjJpnTS81jhL3qNjMO5xAY9sr
Lw7B9Eh7UYSReIrRsQZYQ9+uUb6TiiyPa9o0IagReSrRU/Z7k2Yn5GXtCKxrZQUlTIhZntHK4c+N
p/nQ+C/iSbJT38yK32O/+EQmgCd0yxEVXUzs9GlXZI41wt5v0QCartfaUOIzYtz4fbI28GZ430/h
dIyrTG9dN1oSOALfz/j5H4iEUOuFONEOZxdJ/ul8LQGhPn4InoMyWmQdLL5AxP+tzC0j/wTCy38Y
tTC/oMt48+LJ2JGFr87NUhVfnADzaZNtpqCac0vklx9oHyl3NDpWt1RWcHpRDwhsnfS8dFCG4ZCT
mSrOLtvHecEPT3VGOXuNzgu/QPSBA2k5UJMjosrVA+QGrz9ciqgRQUJr4E13WZIfMCMFkeC92o3J
gganXeQd06T9aoIW22loDoZ3oZZ2JYlrDJQiCRcNn362//sRDOtg2j6bAw2UodJAFuuXUGpY/zGv
7D5rZYak7+3aynkNfWV1yexJh2NN53GW9RFwBCI+kCOoIh3rbUMhpCKZStR3qWWvGSTd2jrDZB6O
V/SPwQ7sfM7IdBV6pGHFP/TYKCnCKVe80OkileyGXNu7AKQcSUmXaVORgO/kIJhw4NyHFTNReKN2
vQkIn+hOt3gnzud7wX1nR7nr6AHIAMhRQTkvENEpfDWh0awH5gnLeZRIUAxATCyEu42vKUmv1zSz
Oh9hoA54s4rKJbMIDJ4Y8j0//2o7k/R+Z0uKP3LaSUj2cAjelaxiLLVhHIrgmjChm2ph3rLLD9vv
zPfmWVjNQXn5JPkguhJjYqNENQd5SKMr7fs5f54vTmsUnHfuPxsHVWKQpAL/+AE8SyAfAIPcx0LL
2jEbpewYildAJRs73ul1vpzMzb9uU/Anvy1YEJceJ9JTnL6zbCyATrXqfqMX2ekf6Gl0VDShFGbz
ECu6dR/JFtmfYr7r01m8O8VAbkeLncU8FIM3XOyR21RKxuOLw0bCOHvB3Z3NGD9jU6VKQII3qn3P
M0g0fqo4gqD6+d/Eed7F+Am6GdYCxkUz/c/k/eP3nVcyiGRhQiITGAB984yaIZdBTzT1QIJh0EiQ
4+XdXY8nO4NIYrDeGyVeAz/1ymZoRoUoc4eSLRmHVJIeX1s/CSh3OJBZAjoRCCJecDJ/R7Bl5ABk
jzKXxizXT0PHWI9Gu+B3iMUIiwjy3CM0cIxsfeeFNgB+pNgynEZPW6QFb0TrMC6PUvoMa3n4kjnC
pHMlNqwRDfNwgo4haW53L3jcC5+zvoqSpLLKxASHgsxCqV3FX/NBbXHZJEg4DJttItAR6/PnDBFx
CNK11YQffGITQrqWE901MJ34imoX4XknZrbrJllg/Y130i8C7ejdAnkPcJdIT6n8tEkwJxHsTO57
Sbkg22TFATRuAhsvEBnnfagi198Ka0u3hks0+R/NqZz8CnwmTGCEniVKTYEG51z9iYDS4gZokkNB
nmzuDXN4l3yR8R8pRsOIXF9CD3lFmjQdm0qx9mD7pGbZWFs7zTiC2DzT9Z2VqPisStkpRB3Duqlf
lq91piM32790EVnWq6DM4u/+dxkqwo8picRzxNfH/VM/kW1Osi1GWKE+dxyD6lRqxgjsFMpvlFdr
NrFveWmFbWE2zagkk5dHhVpqWJb2xWipDIk+hJr+E5iEb3U4Y2csIZ1RJjoqM8vuUUIgLllP/O8Q
0+MIlfS2fG8Z2QYb8A0TvMjbu0q7dv4WHmlDt5HyFvw916mJ5MxKXU5oVO62pHQB/kJ7RMSZc5Hf
05Ztv7sI30c/+eue7EglcOrrIBqZtfvxeaomyWl6YitwU1VKPSI3z3p/dbc1gMDfcr15iqwNCGlp
dgw5eu0hSZ1j1dKSmT86YZSkXBjDkl4aJh/zm9goal28YW315xIsSc2oKiKdhFjT5IUVPlvdFFIh
4b+PZgoRxbWiO21/ZghdQ/+Z5X6TDovPHUEFfHWCuPSSuucEnecWE0Zw6Xotu7CBLqVXA5Ys875y
tNZ7p4POi/qXg/DPRU3Xnwe/QRx/tvxGVNq04C2SUA/dPrJ1oeDdmyK7Kk2R4mwH+2cDUvbcRxRd
I31SLsCfgBA5poDArq1xW7ekMFEowZVdVmuZ7IzdmoE4NjxlFpgPC1zO1XoYE4w+dM2aTZQVRb/B
mnf/mWi968AfIAKec+vmP23yBdamDLeAepICeDfrWRHjBXdN38mjSSmgwuS79Wsk3EH0XEG/BZ9r
UygsaCCQV8AeriuCmVqZbewsvRSbzMKXAxkSi/AXKw3Oh01psXpqZCSNsQU2suuPDAV2CKzIsqeO
kR4/anG8PLgdnm18cLA6DZPKD0X+eEQrBgMRbT2FXLVvNldV8zlAzAIdb0wRD6/xDpOqFAuOHQtK
Qfcu76GUPXkRlFv4vBBV8dHuEIjyLQZCk8iLV3LzD4/IkVQQRdeONG/HyXMsc5WolD/b8MXD/91r
RB0ewvx9iWaBTzlMjOyrqu+yUmbPloO7tUpQAcU6Ws4I1MhhN31t3IwxLymyYgnTecHkrdQDdB72
3I07f6/uxG6tjxh3Ybv228mtwwMqOHmCH99wgrjqD/x+ug6oHnOFYtc8Ofc1uaP4Kj2bTn14ZcUf
8S1OlpTEuFtO+nmTPX+i9tNEAFQeVRVDNCgGl3aLZW/6bJt8lNqc/DDwRu8xM8yD7/1fgc93tUIk
tbFCJrixxeTE7vTck/42gOAk8/XzHtMnWZ1Ot85V5XO7TvkGa0GywrbUB1hDI+TCk0eB7Z/nxUNk
XKM/hobt/uQV96RLNF2UzvykrhlOF+ODC+fh63wdu7NSsdpmuclqQQ5+twZ3UOge9HXIGBTysC8o
onSjKVKVYZIn/dz9jDdaVHMdukpRENPQE9UmHW9JcLILQLAoWEQbObDRY/9fzoJ8Mhx4gUfFmlY3
qbzGt2QQMUqAZJ7C3qRZuQoXH84Sy4DF0KsYLPtuwF9pUfpFh1R2Plt6yfGi1/RvBvweMnD+06wG
VAYyEEgkSe1JgKp4BQQUuH6BcrYCfj/iaBCS4TLsIaYBHv+Kv49CyvMoLtkRpXElfim7FQxlED6N
uZl5bOkPO/k1s6i92SHqgSHpMsmLKguPvqvd9KxyEfflhMkkvIpxc3cnFI2M8Brx2vFkdVZ42HRf
bvsgBvfR4YxfGdL3MtfAs6UFaVrnntd/r4+XJ2t/7s3dg2nRVIwKpNTVfXR5Fo4c/n5W+GTWr3L0
DkbnAvbaW0gF/pvshbq/Vnobh2hokMtNtlBhpVquvt5EuS1R5ZTQy8rXyhYpZS5CdcFjg1DovvLk
YcvMFBWfqaIrPTdGXgRK1l0ACgnEgQgLc/y2Rf54tBx00PgLIDJsdxNpsaRvbisS/6IfrwkQubPy
aEXXoguoiwtxK9s/OGDQZbgWJokM5+cyXIwMC8dnLKMW/trFCkpczz8jfktDk+pMErkUsAQ1kG//
toycJ1KucCeIjQiTSftMj4J2QKXHobgONsfoT1lY/UhFRnNcF/qpqsK4RyoziadwzVGlkfWiGA+5
IScERUUplyaIO5Mgn7jv8NIkdiU8+/CUr2MaPOvIw9xZEipuoAWdHvUzJ0EVRcmQldBMD4mCAjD5
zG9w+7TfCZzEnU29lO9QlvwVqQgrEG5TzwH0r2eK/beNpwjoRrZKc4krkLx44Sd5ZeE86WtjHe1q
PN451JTgXuIXLUtNIUUsgIIsm1lYM3vjKO8FzeoU8DKG84Ti2S1lLpjaTe5F7a7hQurEEYAkkaum
90qQHnH4RfyGohHACY19C4FCSaDC9MZNSrmevcTN/cSLdRJt14DRE9dafTJibjyh9x4ZzfCIl0zT
QYL58VkY9oNRLHqs7Xfk6XFBQhpR/48hinhbUQc0TqhdsYVNAn8AVCmLopJB+B7vKp0OELNTGRYI
sxKhueiqjVqf8zMH/yoUPFKhXBQGfVj3SNjFsH4RDDzGmuGoLNK6lPnl4rFULpLl9qRSHMBS2TTQ
jzFSd+brnQH/cp9bYo0MWF99Z2q1A+pEjkV9jLdzUh1sH139LMM+FoYCOu/ta47RUzEvSn8Eg53I
MbVgvoRHcyaXfVE7li9kTWx/G/HKRuMPDmZhuymuhA9NR8hrGAWh7TEWcoKOIzUhytuqJE+sxxLc
yPhsfyvOTOKuVF7L2NyNIWurlmafgDC+ThM6ReDDEnj4YPUzXAW0MY14L3b7eUGFouhM27e1qp1M
yHwcpw3fbscf7k7Jogy9RP9mTn1zFlVRHQPiHjmLZQoyi5exfpBVDMvpuALsKlo6TtuOUtE2oA05
7eMWaUwwxqk/Wn8RMdfL2lvTkj1gFaI4pY3wlhE/WJ1NB9p3az0t58BVwWlQE4FcGj2X/PGOfIIF
8VL8cPEPOluN4/uhj2Zf7GXl3IMLgnH5YD/gawJX7a2p/tg4tyGjvX1xv1CzX6tr++YFR//Vr7io
A7JM1IkEK38S/g042POfl0BLJFUtJu5e5CN+egK/w4aamI2rjBzpqWA+UWw+qzFKlSUZQM+p91SX
iFiylH0Wc32Ms8IZpF0s8tHbavzy/U+fNx4I8jj66cs+T2knNKIxvJ/AiYK3ZDSCUtQuTKaaQBb2
bLeqwNW8bs9vZDEC59Fp5SMszIwQZj00XzbEyClAoRNjT9KG8EOQV1ehMPeXM/aQ5EuKfeZmXRSd
05ViZm5ojxSP4FR7ug9G+Y+RdKTBwpx3Ahxgtsx7l52Go+Y/DJv+5Zt+QOaxL5PKv608xvWnwpn0
TcnZM9BN+KdQsVNda4oXxS0KN+tZWqDMeK1FilhJLZteHBf+9HdDdemz28RwwIFP+SUv0tec/Bwh
b9Ykd0R5ZKHP+Ikw8Gx/yPBsFkQDhUJY5k/x9q4aEM0Ue2R6xGhWVt29uEgHHJL9TzFu6Vc+Xoug
lU43kW+lA8NN6j5w5Jhg4roiTkEgabRYRQJ46nId9Pl48epizIN73IP0DHrdcONpZRUDJdABCIFZ
Cdy5zQ6OZBZdH5Es7Iw+hSTOI5yeuuBG7ZWD0oxV5hx0MDCMGWo0vSpOA9NNCs0KEZimuaoyQe9j
2gfLWz+X8OQ2PEZ/v01tdw1uGTog2ZxF/Ezh/e8kQNVLX48Do6SkNZWNXR2yMl/xnmmoZCnLBud1
VFnG8AO/xyIoJPULFFDaiYocGfwPxWo+q31OPjMWqNNjcBh22HYJnfqAcfM5ce99Q81VcH+bDjxL
fe/8vanRSsCdtfkdQRmov5QPWwqKAAP3w5wynVb5uY8jcU/tMPXUGW/5SVOnKCgch2c4bRdSgXc6
GZ7msrrq6Zrs6StgUm7cZT1vpHAHwsdj4jnRrI5rkAeNn19YkFfwfpATmVDjHzAiJuGSpqOoaGX6
AK8vBpDRaWIySiHgvMXQPSRH+2XES81qyJ7+AO3LtBfWjBvwU6Xf2uZbpRfcRHQ632TqHroXEyWG
pv7g9RIybas7rT+kpKxhRJCVTU/m7srqsEKYsCzaH+nehxMAhvT0kS2CZF+d0W6BFyhEsCZQxiVg
JC4Njy9ULWAg4xA+6NAXEIGsjB+7avtwUkIc35LRPxteDvQbSgP0mKM4UIkpg+feDGfbrtepeNZO
16IbmsiI2g0/PmycUIeu3MRFVgf8B99WQxCEIGvQqngVRfULdn+nc+UfxKVJVo74X6DOHy6qOBil
88n+3GE1Svt7t/XqB4fp8F/N/HGPq9mS6evu4P/dBTH5J7TeDJlB3ZvE3C4L0OyTMrJKjBFlhZUN
rh2LhM/ELPULnpfMxT8E7jiMZSfobapFr2TzCE4KSm0207yu+rK2ZYkDqzgRni6riqfH7byasmn7
9h2n5gsYylGJj/1qGomMaV3vDYTjVx7GJlqvpxleFrHKk4R3q5eqaB0BSeUp+1xrq2wgBX2c7myA
0tf2E1MAJ14CT+XOm0imRB4r+ga24Dq1Uhncr5cp7Le44lK1IsPQmCEShne57QZzcdeNBjXXFPJh
sJtx//YRi7p2uYmYVNmooljWcMogP0v1QUZWy3VZP/V2nDVC3XCdADpnpmDseCzNma0i3Mh07Uku
CJvm6K6iKpJ4t53Cbx9okNq2UUYUyr1pQ0mwhiDAtGBruWh0LwUYd2jLV4CVksPxpr0nA6F5AWS5
UE0zKEFmcxpEDBaeiTx8Ial8gJyJrQt2jMPwIK99BJt9c1XnS8fj5p1VVRmzazGaXXDV6sLEYkkU
3vC0DfRWG2vNvPTUerytdqvM0RoHTwU694qbfpaG3WgKfZiqk7lJQzxg+dzDBoG8H8q/at5fhDCp
CHUz/QtuX2ofMK0IsjhkxYSl5X3JZBcFw7fJ15PfRIoR77PoqEv5TvZUoeufvcbvtuT91eSxf84u
8HTdxhAAUJu+CPrnQUllTjKsLI2sIOYvgVspa+RIiOgIFdcOLXSiAVTYrDHEpAy+fazxqh5XSE8d
dCsd1XFk+sG/1rrSFCmMXKyg1cF8lkAtcrw2RXJ4JExeZFD+qPgtzKiy3RBjlIsqWiqrmMqdYIoC
EXqaeCBI8stBBaq+2yscJjH3xwWO4NGIHAeme9hA4skDX1VUy2pHuKIG+dXTRLxs503JvS2vXAb0
06+Kp1Zrno94eXFfQMaH7y45JzhW7fswnvbOQu4vv/2AD7GxV8UqMZypV4e0KBaxdf0McsKdC0W5
f6CWzAZ9oeUOmtaaUGGTNXyGktzxEcjfmRNvYE8vs5JnHvdvZ3aCjwbwJ6WMv3Sde7C4TzmWxwwK
csRHJ7bCFqxhfFuNlDZViIqcExTFw44NYgZp2ucpUCh2r4//Ct5SUG5VHQgMwxXY5SBdF/SMKLGF
BwBDO/FqZsxFG/38h+6AdqN2SPjBvED3HCXj/7GeYxfbYXAQ+Z2shyUPacRV3hXERdWiXAjJpVUm
38VrpLY2vG83JwLe1Jt01NnPqX/i1UOvwYoT8eoXxipGkTMN+xpC7aTZUeLSo0CWQgCETBxaxEPI
IvekU62R3YzgzC1lQ14PgorUartfeIBUNvXNywYd9D6yC55TbwAul1UiJhksgJ1kOoiGsog7FlSK
Du2skXFZvu8jjx18Yhc+Em7MTZ7UtPR6Ynzirl4UD9GK87jxj4Rjp29KC/LbtpJ3RCjwKICNjwTl
wEKpBz2c+mP0JK1wnwxEx77McsO7plRZmv6hTx2tPfdFBjNBJt7/rUrc7veNHMxaKBjjS3ZOyyPQ
xw/8PB0wU23JpP+yTV5TDy85aPuuG/aiCLX+jq2f2Y46BOaBo4c9XxSbQXFiBz0lgSi++4A2Vkj4
CzxrURFtFxqAmwF6jazEei7aSUVJ/vGZwm3JdD/Svx4de4DP2RL8Nezsr5ZtQAsP0H6W8IclP6pk
ZjMed2tFDI1/xw4+LR9BKYPum1kRLlR2nxDcW62L1lmrrIZDAQbaOMyX4xh3evm642LgqwBQESV5
gxKf+VKKUGpLSxbRe9pPWOYeepXBAvDPIXfz7fmh2Oqtw8N7RHJa4qXc2hKZ+0C/3+cjn5FjY34p
/kKNYPHWPDYjhyXvp66HKi750OtqKQBmxGH/3Bui7dPq6Y3Kk7nL4PnUEG+ME2f9Nn27STHS9uI1
b54dDZUHpiiiVjj2xqr8HaSbMBuD9Q+eM4uGzYP20/kYYm6NVUnt2YjG99B2hph+WW9yjKEK8ZYv
yVdzdgA5nBlr2IFrsX/yYFdgYZor9L2GdssRAllQv2sgK+Nx69iwJu/FkglMKhfuqppK0uH1t8by
IO3erQ/IIsoCsdP9nxtkRbE3BrwJ/rhh7DUGf/Q2f6h7FL3711MdV9QbkqzVqvDvFeYDZTZgx93O
yM25Hk9MBbzwokvmNwoe0HDbN1ON1Xbco/hQk0vMQnnshzj9dwSaftbkUon7Z9ofm7jqfZEHc1DO
wWY73KOXnXika2qw/Pev6e1DcWOidQ3urKyTzUPOP+gkSCdiDoMnNmvWxYOfkm+JZjVhYJWTbQI7
RH9e18nYVCqVtuO1XkwUrdBTG0VAGOWpWdTClcdUwwA8ugtR8wfsVlzXTyqdp3goSc5wp2KyQOCv
ChZVm18yD5TCD5JjYcStIbhKUo6HDuFlc2n2e8S13p8z2haUSWs7Ijy8VHJfUYyvFcKIhrsbrAlx
2OnBMadHxVpTgeyUzlWpAdaKOGjmcXME4ob4YjJvU5encAH4CTskmjj1RzAg2YRPmx5y/IxIAof/
TcJzM5BDG6hl3rCmEk3YLDlMo4+pG39Aj+V6ugZYXbIHDBV+8jMN07ybKYG94uo1rVa7JR02EFZn
5yJFAFyw5g2fVTcy8pw6aPbyWSnM/b/3Kr/UnJBwyy3UfmoggKM9j+lAGFRcVg2V9swW7C9WoxX/
WiSMwJkmf8p5JGKlze4JzAgcFNtpE1itODPO8/+91UzIOGqivmWvj9wC+aZyukn4gMiGSf646uyE
8qbdcyjrV0zMAmOT3UVFjoWVv06tp3qcMKB2t73MVOUb4PcStnL6510jabw2bwc0A7jerjmP0R75
DQUVbnKmwQMou4s0cA1dNstMa8Ni0fwUoHqxE32GAJld1krfmWnfiMnnrg2rQseXX1vijxcLyyKw
WAfKenIMl1OAKDDXoq8Lwd7lVbLVUT6a0VqkzOlH37psMRIGzcUfy61IzCPNVqTGcw7NLlXSFG42
eSkBZ2necVDnI6Jag0Hc2q+OQ/bkDz6az0VFMDSSPOPgRvwudB0TNDe1B3me5y54WcJ7iUvDLs+U
DmPF3Ps955tLDSyYsYnTGeMUonZ6uH9ZXkKVHf3yxqLJLPLy9KUbmii1t0NemXTg1cSkrDlA2hvb
t2HuiiOX7CksGqUYg2fiT1oUHtGVwyG1ljrwAGhsH1XtiOCe7yVwXSXOvIAOxPNsxHxF+FLT0YGL
XlynKKpNYjbSToacIZjqdWE1rGqVGaBxj1Zp96KdzlIhk1Ks/iw56tDn3dhG17Cz6uifrpVvFk3R
xd5mqf/dC4asVTa+vZLLKohaikJuxu+sV+N6TYVVrm3rC8xaOlKMe2dg/bzYQ2f+cwdLFX27ucn6
guJRuwD7Yonx0lts9LMaNQ91YcwCyCj//jb3J6OAEYvABaR/HQ+SEVmtEOSs9/k64iRMlylub5A4
pKnJhNpnXkk3wjh2+EFTDiHjo2uTxiLeL+bsUyBOOAVx+NLLYDhXlOcEz2dvS2LqjkOBHTuH5eO3
+BGCvHlQTQmmP4CtxXchjamfHFHHNLuy8oc23rElkb2O/c6GfMdk6rAFcDpwjNHiUHGJMP8ZyH2O
pCPF6h6pF4nYHb/9QtyeVJxCRMChSuJPcXT00+Dc220i0Wum6v1VI6L0IZ5dOP2qeASZfDfyO1dz
mcDGyxyFIrkSaCahkWUM8DgGBZSG2Eb1uAcikqM9XxnfF0JyJaz5lmGmO7jyg+YTCCaXBvppe8IA
0sm84ZVtzJlIpyRJrz2/hwKdGz1e1MmjEnwYxHYozkMH5/cN70MKx/iEhtRcTPvlJHJC+sxQUNMU
8JVIuGn+StG6I3pH2voHdG6smC2UciiCm72s+a8VDvHC8Y/7nfxm7dBDSWAXCXioYbYE3APehWUE
o4ux/bjA6+IRsgFPmbFxDMQSrv9WbuBbp5GSWi+8hissmuvnhcRSnPT62NniZ3KdiZ2pvGqI+DzL
Pjn5Otij6wb958vK63EXIxyAADfr3UlCuaL//1sDf/G2oZx8RvbVvsQX+UquHfyIZ1bFs7IdTYS/
8fEzVSu2l9aUdZrM1hMrGO8vnyQ50jMLrso6D/61KYBrpW/iqjj6w1Poc6Kee9S6vycbifTXPJ6n
NDQZ3kDpF01grJ8fUGQ+T9VjCjQzqko4IvvmG/EEdXkCrwu24FP8/9Yz2WFSZD7pgpOe5DQxc/Ym
5HTzXtKhLXJSw42I8mIobTN23vJKJnobi2V0qTlHPjBOUBSlIjZyUj9P8XYh7o7FHKS1YFn6uA1q
xZtcaQHyY5Nh+nID15ey2EKJAj/kn3WbN2RYcEeSXhbEC8P4KQQKOZiVX8VFTBq/K8X/UAffFdH7
ZF3KrjuT6k2XAHmwRo15mMVHJowJ/uswUkTmz9K/rN/X+ZM32emhgAv95fnOijiJkMP7dpJw4EGs
9AMog1GnYzBsl7B/FRNidNb0RGEmViublfQiTEKpeA3x9Q8AclVNrju0WeQ+PE5/2lizHhCF/P5y
5ghluvfLrGAkAb/VCqqdBgMiRIUDc9E5/lTskj37dPtKWDvDbBiSjvp00N8sCRWqhiuQJAE1nHW4
4bB0B2x9OTAZ1NhEjy+hgLfdW7CnPkn6IvbLqfnLMIDQ/XJwcHuWcS908+My1jQEsFH69qRtBUW5
aVPSYjjHxwn5lzTcKoNjrPu56ltwJGHNOIp/jMr29AKnDGIpF1DBSzgMA6MfoVFESHVhFIK7IUvX
D4X6YD6RRwKoN++trQclIMHpwS/a9nDAcPaAckYaUeq5E5BR3f9vU3ohunK7Bzd11yJJoxkBbvPu
XdkL921O4DDLErURNS2mpXJ40He8K7d/x3S85G5zlqp+m+ppiKf+xKS0YqxQktB9CF8KX4kblUvn
2yNlEi2c2FI5P69ydMQFzfJp6kgOGEu9wA1SLAF00mfWQoxWsTWII1DisUqxUHxE6g4BYsNvPA7v
2u0OLLYBrSLq6aMJqr7JJHwHIuEWFHHABx1wcPT3sZuv4QIQvz9I/t196OPJpk1AVVVmEsiSQaVq
Kv8OifEBftGCd06qNj/OatGSDA6P+/T6gwzy9ijOD+Bjbw69Z4+o6ETs9PXQ5UMP4J6jhRZilbUT
FO8H8jpuWtGiFco3vrq2LEAa3+stXCsWeRhrwj7OM2G/WfpVq/lNwv4Cj4/wijMFJniLYuBE3Dxv
AXO/BA7wEjEMwWPwPV26nYsucRz/R4UJ0ISnl5m27pMWdpWKNWIXkpvHQN6sFOYiGEGyON5WVFo3
3sRLLXDO98Hj/XqOHRKVdKNWtAkufojvjsKyassPmHcXwKbfg7vedtA+isf089bp9UYfNPsRxLzT
xdrHou28QExNJQRqMUPRVF8LYDGCxUv35rcXUl4RibWlWNL0esmzSEw3oAZjkpCgX1amaGIIxax5
+pV9swxowd35gru4+61Y62BOG6RrJeLTKwVI/bcADYFjJjsCpNfNXjJdUqEJunakfYlbNZoMMAkq
7B2Bg1OQlc6wUabZZzjTvh2PUfNV8CBvva+bX3I4w4luIJuyvFr4jtv9S9l0VEOiHidfpKkrJ0B/
KW3hwxdrPTatojWhJY97pIaIcnA4SAYhGmoKBvwL3KsQOiyPrf9aeVQBNZC9+f1kEsg0odBZsiP3
CfqbinzFClkTb8sMCMXTWQGbnhHtq0f4pIloNsytiTgTlRchrbatSbsJ6RPrPBV5I3bkDf87BVwj
Xq7VRT8cyB29P+ZJuhMEOPAa6oAtUP4RLJzzoiyGLqMF6BNpIuW8VQPVStwozHgL3cGnuBBbfbc6
6nyfcbZW7jW40+5341nKomQpZleoea8Zxd+Gdg7y+IfEntsJIYeZ9OZ5MSHti0odXQV+bSuP5M58
6f+pv9/h7cvhuFtvjWHCxkvN4g4Rt35FomtUi68C5Z+MDl6jm705PTV6ZoqQOVEY51ir1aWKyR3r
TA/3VET2ErmDDV8ed1/yC8E3QVEKOXsZWhwyRgbGCK1ZFMEeLvHJiFO59ZQwsWGo4YqkprixvZOV
zw1UWt06xRQCPSp1LPUeUUcpTFe8t59mZmG6GmNWhUDWsyuqBpw45AakIz7rwYfxcB9dbQUtOYjS
1R8XfDH2nM6t3G17ZAvfRQZm81k3PlxXZFcVrblko/ZBAaKRYiIECdoNt7xUSL+bH93emgxRNOMV
UzA0CX8AreJDAW6nQwho5a91aCdSHL43barJNQ8RgMGJj+UPl8ho3CtL91k3KSqHbgENKmAPxFbe
J99hM8+AqJ4eOq0BDGx5QUB220cYUPfQX0GSnRU91Le4ElrtXRSVqBkbSk8Nolc+ofrHked/KqDM
JlFKk0jGTCGgFVckDgeM5kG7FhKsYm6kTtvUIW/mvSMgr8MkGBMXY1P/cMfMcCQa8alhScb1lVvd
nkPIIdQS/eTiNJuykudhBvyonJF59XPj2j+VRGHzWxuXS22P4IjSvAJ6Im0rNqHmPwJ7PizG14+z
S1kMEL/0uttxAXC2Kor0CpjJLCAdfYdyUu7ZPdy1Unw7WuOnp3QiSs2Xxu8MQiLwRK9Jy2ZMM544
KBhIu+GnfGXZizOIoaaaYqcLcCJA4aYcwlSf5If1F/0AExyOdzGpXvue0fh6o68YrkcG8YgvDxzK
d2wWfNfNnvPkkHbVs/UpGX1ya+yvayn6QEvwJLSbNjIAjzyjjzLf/D6081fT/fefLXUAWAjPLQRi
s2U3C7DcYntOJIPfNWh9Xoqs8kJfVeH+5weVIuFLymxirUJO0rHDbsz3bk3V1eg5BdodmLi7rAIj
iHYpyQPh7UHoCoOAOwCmDN6RYyKMKy158LgxCT+HFfNpNTvwzoUCmavc+0UhPP8Scg5dqZM8IoEj
9n54JUAEWWmdEqA+UJuW9KklFtxUkSAT5HSERypdkBMh+S8VgMmy5499W7WRcAV+oZlCArZBDsvm
SF0fHODJ4One5ihLb9KNog0B7N7sMbLf/VxK6QAoLO56A+HSSVc3OVyaLBo0w/qtAnMwuHOPf94q
QrUyQF3iskbwhINAabRkPB3++/yYbli9r/Xg7c5j5+X+pES7Hz41sA68dWcWM78k2W22ItWdu6Ug
ddkwjlnu4I8/NQ6ALNayvBLF6IVduzBkwFMCcXdxWZdJW4zJWQDcQe/cMb0USExZK3DKcHHzMrYt
Tgol7QKHxHC4AqgggoRO4tcc2aU3TtsUBkfYL8mKliZO4FUGssGdyL8nu1yd254vtSKG5QxJ9nhQ
rsBiIQD2WtR96ThA/lheFxSu7iIW/4Ga/ePVLmMiPSlEMdPnFW5fXI9irWchiqfmUFbZHxu36iCK
boS927Qqly5vQ6YfoXRpElAGZS8xMYptp0Idq+9rlWwBpSVwB65BX2w3tDt6YADAXUOdVf+KvQFl
1FlmEI1CiqF0U/sV7qkE/6fpmr1ZGI6ZxN1981Gry28orf2jsxR1B7o2DPJpet0LGfsal/DZFf8T
eIb0iNFjBXbg6lV6HJ4PsjAKTUtvty0R8RR4PgCQxOnSmbP+esqXTzr21wYfuqzpU14Puii8NZLN
3jm3bVDQlf5oe/0fqFsz77hPhNW8zd68E1O2yEmw0NWgS0GWVvYLvAk2ZYY6n+LKwwuT/OiPTO/q
x/UdKMshrHuKPxWHJx0Pth8Ai+uITz8vFOF9h5a+FTrPZq5exfWXS0EAeCk6DxQFXllJ+0GRXGwp
A6UowjzZ0Mdoe3Uloz0xEyKeECp8Slrw//jobEsR68dAvnscNb/62c0V5ve4ixG1DCoKkF+VBc3J
bWZDdFf/gQVq7Hekh1KuGwQwhRJlmGwYxhF4hZxt0jjx5ko8sOIWwTmzxuQWJogYlRNn4k32YG9S
MbOOQCsqcGfrgjPCDDovvOS7J9TKSwL6T8TLyHh5BL07b+ajEdOX/azIREld9z7vl/uBVqcLNvcr
hAEbua3HPftlRCG3Ygsgbcy4k+W0BIjTESFLs/Hcrkpu+ctwiEpRYsXOGMalBGNPT7+9tZgESkV+
DvtPt0ityXWaBYQZXTtCFiXOFH3p1eqT1W2Rn7XwxC1+Z2g/9QmaktfBcLXqGAsoW4o4jcIs/9vQ
vtoYzNtlUEpGcsmo4JFFQ9fwkZlJZ7lHzScTBIoMPv8pcY/Dg7agKUycCxNumbkdTRkBw872UXc3
IF/q+9OWVJXZu2rxL2zgK6kA4Wm9t/K0S5reiun4Qe/UlEXO2ELhk/HaQ5xWn+WSB/DLn6+1KsPb
qezGdutG6l9892jM519NrbV6RhzLgbQLC58hdqkEEp3PAiIf+tLcISUaTdtjDiljsHRko6HiMScq
OHdi3xZOkQEegAogy3YFaHnBKYL8144NWcq4MQ26UtTUdUXpZaN9bcXK3Kn9QlVZm04OflDnwkB9
z5N9sIDht8oDRJKEkyHQZZqOIxJyQ2Pz4PSTWBWHvspvxyweJ2PR43G9Y+/D2phyPQpBMMZ1pPpF
MsnRocUV+Fkl2rWXBzwZt9Gjgsy3IOnk0sDC5ppF9sC3/y5bYh8IePZ0w/hQ3CT5U8PHJg6AYoV9
L/eMQT3hTo+3vloj5jnW8tbyuHIyYUECiI84aAt+ulV82r4wfkzFnC8ul8k3LwgcKhMfsvtJPCTk
cjkwCNQo9cqGvVRtCohQbQDub4eWfrxuRg1Ca+6T83qkAnRqCvyXcN+I42c7E8YkslXE9rPcObF0
RFpdR4l9GdWYR8jiLD9auPYivgQwVIUxnr3OoOh0W6XafmU+5Kd/S71tUhvB4I8AmRPDoMUAyddn
Msj9KIfKbR0/+OjXDW3ugoYDBIycmDUWZ8uWszwVhSDtmnF4c8Ps0ShkS+5qoBlS+9phS/kq1EDB
jD3kV+S/EWWt0w1Sm9rgW7Imas6QDbO6aWXtN3ZdWXu7IXjrH9d/hVb1FYX9WT/bfpuOdASbVaC+
ZrCxS+lfxJulqFQrT4Gwysyq4GSkLtoaQgQe4hIA7Apc9ShtxYxwtU/3RQcUltXjD50zchMkcSps
qmArGGk1dUy38qHXYS5KqoUj8oHj6bRbMS4vqjY9mS/vQAoUiFW3jDzikftB7DRlKaUG56HEqn6W
M5C68+9xn0RB3HzGaYApwz1QWSSXQkKw1qf87Z77iL/9uOJLw0MOQ8T29wNtQtPEyWy2iKjb8u8Y
FDSURhaqKyybivNKD7vxAPH4CJa4JFwUiZiVOH8pdvuXKhKrM/dIu6lDexDw0ue8uGPY0/i3sxox
l2VaSXTuDhbfwzKCeHR+8naQzcsYUPT8Skh3ZRv+WGiCvcph75gl2shb8RW1cN3eEtHswEgrt6Fl
kuRRZOUpATU4Tki/Qz7OBB1olBLjY0jlLFEdtGdntfa5jcJWBIdAygcNrRC+ST46IWC+1nZXOLh5
p/fSVLMDwt+tsokx8AToOU3MM7kedvtBo7PRLp+Jgopuova5Gjio46NvzdzMikTQQ80CSniCXMMl
PnDx5CMZtCMjHaA7ePnxbEYVF1nvCpvgOPNZRSOkVGpRT73rxSHAveghkUsgMfF6d/BHO0maoIwj
/77jAPFAr/k3HlvjLrg7wDCTNuYLlOUI9+TyGb7krGzig3wAeqJBcVnq1no9E4d056dt7enFSW3u
w4XFBCDcBpNyVBpbXX1xCYWr+Mj2uYOic0oT/njM2UwCGlhrJDQ6mRpJ3AAT+CwmHcqYlkh1fDFB
Yt1XyqYDK9KyNhYOJt//8bkdwAVJhd+XPoxvCKKDSzawGGY6bItvpbhFB16mhqZxcNtsv039hQse
dH18E6fsZ43rUmGB60hk0/s5ocsNM51MAtvlRsZ//BNnBlFw7lXGSrxKszsd4HHJ9rQhuwrUPHBC
oyIsiBn3UiB7Ohg0I+eIruvtu3WppRe8ln7lAE1oP/QVqyvdr0d/2p8X5zdMba7/+Lh2JyeQBURP
bN3spY4kp8Q6xaehT1msxdiIUrnWuGGQ5md2S9RjUdNfIACVqkndiqCFDzV8++9m0tz6HQbbI2AW
XyW9PuxFsyivvGwVtPpklBaz82q483a2mX+ii/foE/R8u1f8mb4Y+zoOmwuy0doO+INS82CJZEMS
MoZOD+m6sWT3CFvpseqPs0L2qXEcwnXANcymSGnscDfj0TifbtDSvY+THosWwptk+JL348GOs+dd
nUW5asQMUhEK24T2TJOD7x4tELISMGHdO3YxHh44kK4JTk2N00KP1gnJu94xvt+0tSUP5mnvMWG0
U6s83Z/YugMFhGld38XTR1MCMSjLuTNTPnZ25+iJKW1S+RBtf05v0rxzygTj/2OIDi+n2GLTTLNe
FxCr5cNoDwz/i+ifqZoglQF6KsoAv7kfo8KymqSx93g07PLI1GDmp+t502PeJAa7vOxmBWS587po
+FLjfAx824KSCI2r6OO8yUEX/ztqMP4O95lLsstU07OlfDBROQIqeOXmKwBjpnF+2EGuO/3udMgx
9HO4VDVVwuyopcVb2oNJ+KyMF5i+g6ytcQSVRuoHPcVc/ulb8CXOGYJM07Hg20hyiOGbJ6zWcFmM
u3G6fOzwk6yv52LWGBSICWIoKB+tFZGefeocmX1Nk4thWRgnNA5kMj3Sv/4atuSrzzpuj5AzmfbM
GJIyttxeNnMn/RNNDP8j5YMK51yAG3UuCMW6qRk53fnUBCngnQqvrmIokovLg0f93o67D0cafXBv
lIX09t9Ep2uH5aCaxXkuK8N8c0P2JB2mWlZs3+4Oy0Ydek2N6kY6vMNVViex/4gFflp8IjZk9zdv
wOQq+qJWmX9NMIHd7UkSI+0L5xxyf6POdNt0FHSyNdYeU8K/35+40xHw3liZZiLvZmolVm69WuLG
julAAfek4c1jRwvcP+ETFfCZX3FJYsnHbFWBArW+W717t8QPyV3MqrumDMI6vhStlwfDSXv9Xxd7
TtfQKwju9fe8lvtefucJWhS8fLQ5fks2wL1zb+oSesDo5DD/PHlAzSHkNSTXJ9KWQ0w2mesrC/IR
4dhu3jrpEKXMLQOFHlEMCc3rC6JTA2VxuUnpLl8MVUTh8D86oLdzO/jLuoWx5tltYEqT2bRC9KRI
FSPcOXT0sBYUci0clAW7R/XvMjpYL7gVwkCbVdvz/i0od+RsR8YtguqEf1QBvG8nFhAu79BeFjlA
UkwmEeU00NsZK+VBpX/DUvlCLpLxBBNcdRDG15UJW7cj69eMxYO/tqgMvlxBxt0Gn5EAKnQoLZfa
u0nImA3D+TayC1ClIGIo+QQG9NAhZmxEBYChMpSQkq0hU3Xkwuxck17c0DMAdvfd9lEghOWsbyrY
An+8k0OTBHGEY0QtE/MSAH0ZFht4zq4jZ2kZthM0TZjUEX+kwPUsbhmTbTDRvWIXwAC+WCCvfzXa
2gIO4QIn6DlArQr5wHWSApcSCwnNU9eZGtAXx+mmfxmeBgeroHVAgdGM4auTXWUP9Sem4iSKj2CG
kpOSUj9NUy8MPnC2QPWVmHYncQwqQUWMZjuIoA/B3bJhwBkCxWx4jK1ybgLiMflUB5mBwNx40QTV
F12pAfcm4CpylFJUqMr3yL3/0fV7YCx/041GvG3g1ZmA4kIZ0x0OGYad4qW7oT9gTqDuJxqf2ALD
wLUFyzG/mytZMNBihoFMpeZWQe6CB8+l3xLf7EtsMJrFy1/qClSQwb4RUyIcEKLqZ9pQJr8qQAxf
HU05/1lDFVqzFYHVruJ588fpCZ7MDRQ8pz32LJxsGNGD0rJjj1DjxZqC5KT+vJrfE8huAiUEVq7j
F1KxLMItPgU7pjfttntFRzxgFDRvlsvRPcCsZGrRxxMXjIuJ0UAc9BprrOqynzGfL9uZj58m5m6y
v0CoE69fR7tQAyjHUt44WngvNjY3aEEAZPM4hSujacQ8HHza0sx45qgjS5PPV9YOJdc7XRZkp+S1
xS2pxj3UMnOdSg/W3UYHp0Sconw8pF23NIKLohzR8O3k+YO0yqpOSBvJOSsRC0ZJVndvCsUeeU1p
eQD3HAy15Io+wgxAMYodl5GRrNfdJzkeFKAxcm/6WqjkR6vOUwUxeV/z1wh20tDYYXDoilocsdFa
rQZpUKrbMBk5OVq96T6viwO6LAIXm2RyOpCiLGkt2FU+h6qw5xPwnLP610kdXPx4Ewqj5lJ4Fpk6
l+rTFnTZ6Wv6WP+01kmtYyZceQxFo5sxHC7s5Q2VY8/5Yn9FnZzhlEsdybWeX+e9ca2z0XyQ93bt
NTZKWdbc+Eka7UsdgnfIZLdU/v5cdoropQgfV7b/cZq0i3hS/OBY/kq6RZMa8e9FjiFUxGzFbl2R
DsNN4rfIYGhx4NDu+kyNoFJ4JrM65ac0DVKoigh5ZptLrTa852aMUmrdI3U0Svp00x3kUpBSoAvl
UoJe/xW6kRiMw1C5RUTXwLql1GIbum+yPakPELwrKf6lZQE8Urq+AZb1SOjLrQInRKsm0TSq53UV
E9wCjtfxYtewwXBBMySnVBR938jnpCJ/nuYUKc0Z0EJDlwZGVxl09ouMXHvV6R4UZp/rMTiPMr4X
Yr4H2djB51tb0xBgvI1J35mmqOQ7gZVrBeR/hRWEH4NyF7bmGRvBjxBXkg6azE60JRaxtzLWscTB
VbGFfFM6ns/RAWQTHhfNoX5LXCpda/eoXkOgv8D2sxiaV0W4bpoxOIp1l1Siq6qP9E+KcXk9d1mt
dr4gkAK00gma6WeoGzkLdcIX38SY0FQMCA//BwmOWgyjV8loHc2CEAyUVA6OpgbYLBnPeQySkF+m
qvAk9wiqq3b+83029vZLSIomRyU4DBmZCzhleQgoWYOZhaFyD8JLeicjHa78oTaKX89hQ/PriJzr
pp+WqV97l3wJE2L2XheViDUJvMvQ6Ynvjoi3ADzzJtHwKLfQTqdd9c3rBsxji6PIslEH5F05IRhI
liUE+tlSirHB/Va4F64Skmx7prTvsV/+fYH7c84pFed4VMpysG7yvg0u2lo3160mYdWhnomJ5fki
WaSr6F8Q/YvvCQhtGuG1+KgxM0QXnejlx5L5Xm8HFp4YgzyZ8CtbLgCzOM2BqiX1nO54135Rvgmr
fjalKbnbRClPuPevWvEfkfEMFZ5rcA6CZqjfIC/YAl1f4I7o9kPZbfeIdZVflsUUiqqCO4vDVsoM
ZGce4RYR5IMbXB+8hG5h+VajIR61VbdzU1fQvsefibn9lRT6tyGOaoSfEtRPTg4HCvafTLlK1IZS
oceBRBawKUh+W9E2MIu5dYCmKTt3RGP9HB/lLOBqKGsRcGO7bbfxLOBxGsurQxvAijA42N17lwbu
WwXUr8TMhPxF7HwtwabJ5F1dwQ5Cp2m82J0oFEgWM9zaGM6bkjYCtEsIrPSBs4wp5NxQE9hwpIEv
grZyyVLjqzt4czVid+F3vNFn4oGSlTnRzQccuEMvZvZKXGHqQCzLLoAUhU4OHFfzfZGFnhf16NGE
IHGq6c7vY1OlEBQtvPuHLS5tpdrDbWFDqRGCR55Nek+/FOxEDKZ6PGIAHuizWntZDBXWsAASbF4R
GZ41oopBNMaaWuAu0kH/cpAI7Zg7+8GEpqt9eyBVVuDxyEmS5+Xc3lDeY1hygU+2MlzIxh1Fuveg
1WJyJ9SmIAFM81TS7zILG59uZGuZx+wTHLmuT3Q4/PxyshTrGfbFv44DResugcm2OmScsx1SRz0Y
0lEs6y8qmnl9UmnxVPcyrhVzrJzkYQVXWKW4iK16MfhDrDKCs+V0o7qODvjcKG5d90BIWI5eP3AO
CPcJXFXH/nZ+TYXkjA1qBi3Kb94I8jfzH7koXPOkyHPcljQZ/vdzvTX1Y7fr0h0WFKOJY780nBv0
iuJPPpN5BjUo5QhTNEwT5kAnnGzFOeLGiuNytfutq99hN0Q70DH/cO9GywGv8XREqgAG9t8vLGhI
N+me5CQbJq/pjw3tzIrZII//TOyxf+fNLCJUNedJImmVLc1YGwWrpyZQQZRSpvmcmuV9E8rcDtr4
Md9jHnZywqEwomd8zmsDW5YwgRTeMkGPVkKt6rMJSaMeaWQeoQv9G34x6RJmxbsKwAov12AN8wT2
szBMeov/8jd80uQjPbwe0Ve0Xy8BPUfhZd9I4XB6f5zKsKvNZ850LzYDNczXNtDVdWTJrQZu2X5J
xRyZnKid5xNqCl/eVUoTKLhJGpKdN3LXJh0+FvfAdU8y1s8VXNP0d3uXtaay0bQe9hvmQTKUBZKj
J9/tTcpUXAgzGSy7/iKFLrszGDNQK4q955E/sSz0RIzFLIlBdosB/PwRa2zcAczAtuszZzs4/aAd
Lzx427z0gK3Sst3Z+WPt2D3k1/T6jU98AZNIIdZIS/4Ky1YKUdg+lDrtmOEBRogXqIAYGYN2gA0x
2lTk7i+3MhKg1yT0zyg+Y8kguNjJyEXVJYtOywwHA61vHiRoPKVYrej0N4FpOfXq8jdl1fwpy0c5
k3x80i5FuAykJm0Ibt2dr5BTzpnOqnZHKVly5istqC25IUSURkLnb9pi3Nq6a0U0DFE6oEfl6/nj
oUbAC1+ZwydM5YrAgkLFDEDCTs6NuXob31nl848zvmrn1I6ry2fGUxNyuG5vl5HY+wE+3zosRQ2h
d4dZXScyocQmf/ZWiR0eH2t+lpUebKD5lYDylWWl1Dg448C44DNfOCxGWVk3NU3yIVRgDWXQObCC
idiU6fp5levY33NCyVQcw2STZAUpLh895jIZaKLAhNdPi14cht9p1nPEOes1NLEUZySM9tSxtv+y
Nr3Ipu1s19pHkm1CKcygwgvZBaMTdhQfBrncqM1NdYsSYyaej+aKC0c54aJ/D4094Jdk4oewrNO+
h9fiL4H1zpw/ENs8txLHaevpxOGNDfMGSzyI7CdECpdmd//ZM6lAGOU2a6utIbidxzL22My/AgpW
32R6MubdPmurVrkQy8tfQHSfhDZ8Fn48pPatlUPkGp1CaE6KLPX/NePRDFcnb6dWENfIAaQRX97t
cDbCJqe7FvNFPv5lNdzCso3vX8arFMiO35hvcXXKmNNwH7R6i1auTVpjmh3UmCR58yvimgsm8UH2
AocNih87smWXb/kxA0iabtY3RPBizDl6aZkTIm7g8PLHllABK21Z1CmIx1oohXguZyIJIfTtftrg
b2FO46VbiucPz6mFfcyECEgxPyGr3bnpBodQfSigh8CbHzc81rPuMGyBTCQMUPEMsvQumubAYNhV
pMeQ11NfeRakFB/JSl44ZU4U0t4qjl4My+kV7m1SGO6BeKTfwzYwK/noT2+e8NnmTOw8OwxFT/Fr
MySApebzimMGgFw9IHrZEGVe14OIfnNUQM0IXEppvE4+HFgcBl6h4FICrFa3cGNvKhb4aaSSJqYT
1Z+cmSCiZiyQco005I+LBYZhjv4HXpIGOAll4HiTjgiwCEaZDZP6ODeDnlp7F/z52SP6b9HOOcu0
hNwO9h01EPVhA1O5yBGiMBTvsqZt6a6eimKwLVl+SgW73DMEzVhvo7JevJ3n+owuwDANx7artrLj
aJUlmZj5QQxNiFa6fvvADo9g2EUFm2PAd1gYLqKMT9+w2JMtQABWPgCiBZyVVFuegYkW3BUT8ww6
zmFGpS/5mz+vLyAURxCMjxohxHWZs4UkxDUv7EdOmWvRRtcNbXdGa5WiGMeCeqfB66/SNakU4dim
Sesm7p7WhnW1UKv6Jw1megtzQg9NWpsDnaRI29V0wc/r9Ur+7QnN5SjH0XicEUcrccWxDSIdFhY0
79oCK/WhublmKMZ8oSvfutQXE0KB2QZWHAiNvmKuogFongGKLQIaiP0vEagdXv5DpjqlWYBvNWmU
j6y7adRMGLAIcOofjJQTPEhHexmxCZ+SazGPsBwb63vlEbY4FRazE1wsCD/RSnOhfkhxAWMYbAIv
xwDujXPTfSMZXQx4XmHYlp+0LYjP5HNfi7NyZzH1S5uH1rM/6mMN9seg3SWeHMVP2oOpD6712ldF
4LlmxgutfMEDq9L+AmeX8tCuXXJ0w+DsQKKexPtzxP7qbsXp86pS7WX1AeqXZt/e1s7f3W916CwD
QVTfssrSg2VecY/QbkX+/VwJwnvZF8dGUO4J6K7tQwgX7pQxbxyYmVww04Tfp6525LvyJPA5OFHf
ZJTMa+xapgJNnBR+vDzDDYLPxFL2aP400iKQVY9FlmUNqW0vfKstHUHgYtl1TSOpMwksRWQ+nZ9n
19/Krkug2fKfZH1gOgJFE4dMRhCePTHOQRGDSs34aRNwRNjVXy+RgGCrKgBXTeGu8zSHyqnpejc+
TmNp1vcdtvTXgX5CG9KLYNwVIqHMtH7sMVbXSZRJyvT8VUyGxdZ9ZiW8MaRQ1blj4A9kFjPp4943
FImE112rw4jvHt5I9qLkgQ4mpOG2IXwRhYjlWEokYZpehH6xAdFZD+cBj+YslEYrh1F04UxIE4jM
hzqh0iOxThC3QdNVHrbdIRVZylenWUWha/2iM8ST/gzIuyXdRrOC0T47Bv9tothNj6yHZ8Wu2yJ7
bOO//9gsNI5minFAFF5E+P/ALnYd3smXRVPFTsUnHH3nPLIqXDM6cfC9hFGJEpMjR8qwzlj+4mXy
p+BtIg5CEEYJ6NJQiallAV4oNCn9Ym2jprnLDbfueZT9XYX4FDpYmwzqrpKWDOFfTKHlEh/pa0iJ
06yebz+b4K8sBwt1Zvbcc90cT56mfPoYaHGVsqxyED9cPjThzHNa+skfxvQdvp9lL9djils7syag
BPWADwk8dOEo4L547FQ9Yt9Q6L52KOQkm+TZGg0SPcmtk70S35AsrUpqlhcMgTQg9fmZEjPgNZOY
+V/WGFVEWfEjZDJqk4JnKzQjsgocTJDcE04Pf+irvxd3cCSxLVuXyYTEmOZkG76inOL1dElQk2nm
OOGGz6zCXdsXxwtmxV13eGaHpDGuEqbuxFHRl2AVlb//SjbspY70F/u4WVZA3UPmgbA9Zu9DCDyY
TwJYBA/0c08aPtsH+ulFULZ3Qtd2S/TdmOhCYj3UgJgv7GJRH9TT76Bty+aGsIqrhOWuvJxpIMtl
vWxK2Z1cOqtTM4OypMUmsKxwvhI4NQU08d+KJd6nGDG+FyjQMdbXoUgudAR6jm39qqY5ybAdG9K/
sFAmF0n6yNHlI8uH/FaOSS+sR9DDP0lhCjcdGPq8Zk1g6F0f/qZwLymhs57MGjnrZCbRlCVE9cfX
7nXt2LXUW3RLqgtiI9B6wxJr2xe2QimKio9A8u34VnMy1lvAyyMVBJHSaEmu/T8sPrYidVG7Jc2u
2A1LNAjWRQZ/trGXJdDxdxOEadSwHjCmi0VOe8dF5Wu8FmoTG2ylTt9cpdP1JppbixSjKulj5NKx
r+P+jJz8Q9Xc1JmHEMjXwuJtFSj7MzJZHYv1m9LaDtdS4CVhxVuv5Mkdtv1upDYRVymOuHfi4WY7
OrpRolK1GOoINy+iRJ1/ZXRS0F55avOqioNsEaLUNZF74B+tLYIER/OkZf0IS15xHrs9+Tr2VT7w
5zPqT+tK+xFVnJsvICvrxPislBcZ3k63ptg9GJQwCPGh/+UpfnlWs4X7nDf1tPMRliOxa74BVF2E
F4NPEBZWJCLJtXv1kXfUpYUx/hxu1QYN9dlAwdg768wTgSZA+NFiJEQHsoYLEkE9PQ23D3vOL1xv
C7UcutirBbm9Rzgmnz4W5Byvr99D+0PKt+ftUnii/wdS1HajapYUOkxGWBxp4fcoP+lVjwyZ+/yV
P3ILPAUVlBYNxrdz7Kb1MIQ8/CZil0EswOhkajZnHKbu9ho9nNsC/98PA4SWGYQUX3CjdA8PLfEA
E7DzlQLL/Qt6UDnuc3wqZL/3uij4K/IYA358ZEVV+iHRbfxdyGjkPxLnhVh8ZunuTiSzBsfaDYjk
XDT3fdCEt1lfwrhzbvrDf0FzI3XkjL83mWnaS3fRnb16jtLj9ov13GuXW3zD5W0lev34P7hNWKp8
PApxuyn8wGd4v2vXNT9OWyyq8b8wx4bUjIxmLGMfTW7MRGeKuCI5OiMhkKCFQRATDTyjuSqT6aHz
bVDYLR+kfeQXDbVib09WayUc0AGTQUlT9+fpfBjGlCDoY5VeuS1C4fQG+/0YlRqLWfi3r6EdnPCm
Puh96KKVPCLuWhCjmekGNd0gDVVOjMHSaQoGj9tXm8ZHI0EmhNosmvSrEhTZ6BJPJOTrJx5W/knD
mmjIm0V+aSseGEmR+pLo6H1U/yzml/XFtBl4B8lzHG9fxugH7SoQcKkWxTnLXDYsrsFjsTm+RPya
ReZ9f64QTREw2TTeFWHOyNK42QbOhl33YPC+TkJ8wZULNcco6iS1F4Llr5cS/2oqhjj4yFhmxd47
EEDilSYZvoyd7+8ghnouEu0BC14wUFdxE1okOL6BPDys2qV4Ksx8ANuCIHZY4zx0erI2Ntmh+nnN
sA3N4Bjqqu8M5q0pcrN1Bzdege9653RWSfNtjf0TzcSJXViO6gRJfXNL4nFGus0zWcLbdvBDmrki
znf3cPHtluqmSn3OWFLSXpI5XRNTJLi/K0FYDF28LkF+AohOUqv5bsIdt/l00LCVcexixdiBlyPx
ny1Qo4l1nbuBZdGY/vFWxpqwaRdkGrSUgXGGzTIzqk6WizffPQ23oOuuotFGvNTo0NfBYOZ4e4BF
r+jaX76h1RstEBfVt2yKCtHixAR5j3LamIzE3UhqVvhIOnvmc8Z/L+6iv4gTE+IC9tqMEkpHPr6q
4okcK8nw71JOCw5l+A9x+Bj3HzkGxSBjgsCe7eDVsU6lOojG8/7rFFeziLybXmJcK6aHu/ltanN5
smrHigaY85EiJLNPunLQWWhu8guv/9okRjSP/mpwniIfBPdgzumvEXy8P4QEQvV3f0AbyY1OAlxj
Q0+DqyVGxDoUe9+JSKBN/NwFyW8WV3A0/77wKLX4/s6QKj318T8auFDsjOZt5JScz0FupcCpF5jt
uyDLaysHnOLDxCp9wYmZu5pLiElPrfsxlSIUVK/jAsSn2H+NyETJe/VK/wEDM03aN+q6yPb2vV3X
Bsv2Z71R3SlUkt3fDKbYC+tVexUQ3LCui/XvKfedwSmlhWplwxALJF69OMTYsgbEra2EaH+RJ9XX
pILHSqNwv6Rc5ew4wS3wDVBbZRR7WCNupqTFXkQr4aE6hVOr+3ztOyFEZ/04vtIx80ayR/C8nXUd
ruhg9ab0P6rfeXe2b3g2aShC511DhVVHrX47qSzHfHIWRwJPY/vpxu6YqfVTObXb+QuNr4JRlPGT
jYP+S0WJ254S/C8L/mTbDg6hvt00vtJ+Xxjqa1orAcVBLZtG9ByzTAIQz9bawTEQII5f8uuBwgfb
2yzZOayu+i3GeB72u55Kc0iGGRZfiMBDX6TdOyHRZyGJcHgi8hOWWQPDd5xKrj+7hxcefz8CsTJz
MsAtNmOhEm7OSiFJvh3CULElJ9Tn6Pcen6XAUz3DqDgwF2guyOwCQPsaA1AlOh1EEChZ4D12L3cR
GwLH1rABh/xdwiMrLwmBxUHFDzEo6bADn0e1vTddyWcnzgHW0/uuGiJSu3TL53mWHNA3YWOX04E7
xRCApnlCMupcHWCLNMe21GNXup2kGHDm+KrfSFU0TkjYcEHjd8yIS/t9PF2mCNHxbUNYmEA4RdQ7
ocPVL5Lwrg6M8HxJd0muzIix/SXqEKHfjcG5B2fnBH5tlyBkw+wqVdDfaZ1YGFvADw+QaG/dlwCi
C7NRu5nkMGEGu5bvJA4U/XjJaxF6HxBpIrD6pJevCprDYXsM6Tyj+oXXSf3Gm8A91BkfjHXw0RaO
j8Vkm+i48f0aQ/P/U75Mje/0K6y3534Uv3tvJ80rETV/GzyhE37ie5HUOkOWZgVFScpYhEuuu8Qz
aBfm5Lg5nFFN52gPNA/1POJ4+NW4VD6CtWOWqpYE2vx48xw0Dg8PFRRP0WXEyfbz1lrx9FQwcobC
BHw+B0YLnTdPlrAesoogCzQk00kNrELF4uQhFF9d1gkavYr4BPblNaecLe6ZhWyrUv/c8Rz88jDA
wspxOWYuSYNFV7L1w4CFktq/VyD27Am1oZK+vTpCw8Q+mxzvMAEL/RKvrge6iuFrlgEjbHHM/FaG
vKqw2rrr9ueOlNfkLEVyaPrXP23XJRAPHkgGnskLKWrAmkD9RLUyqU77uyw6DqUOyaN3R4h90s9L
LPaQZ5brOMNXny/etXQERxX+mfsi7lM/+n8yZQNVvYsHEULKn1oC7gb7KvUNLhq8tEPIRGQi3edj
KSnroMOKJ3+CFbfR8DEflI8BGEAAJ/V9PIaOwKJPyl2i5Fbe/n5XGaFQif5pLMnrcsXEXHKiQLmW
i6XVu/oX3GhMdA3sgtv9YNDxB+dZU8bR8YXnmtqkStJcUuxjgq5MOs/ZOYw9KgrYkmIOhbx8142F
5H/dqIr96gW4VDZHfu5I968vG309CVKcqrToI/SjGsLgaFxzA45knNYEX346S8/iB+jWRxw/DdyO
M+eUDrv8otDc7KNnrCTj4yvwEITCNCwBeUz6lUFT2vik/RU0bKPDsE4LB32AUkjzuGe8xqEISV7i
3hvKloLa9jFWO6dnsCoHUAvsNoWfIGNXBL40/HPZ0MJnlNECbQ0zxUi7AykWDJOJitvy2z/xehtD
FjMcyJsAp7fdsRb/huwgwkkdeVnz7Fyg2VulT/3m1zaiJVu8YUZRymJTHnm4bfepv/EFgtwk5aa1
NGFTHBAHpUmsBnJL8WgTV9QLPdzqE8Y0PWjeerymVR/DJ3WVRcyFkB5o3nBfQE5xqateSF1zOiuA
XQybt7RDyxjkyU+d6h02l12IlOHq3WkvnzIBrxNtOdee3j0ywu5GNfoan+G4CRfeEPRTyYniPRkk
iheRLSRcpXOh2EYxjBIro/YlxMZ6evXayLjV0lbVUJNzrFMAAi1V9vX2Rd3XUjUCh2i+abk+ptRs
wHJkKvqvumzIJ3O0Z44sqw3izZ01WgK11IivAhUB6ySFBGpFZhCXqbY8Ag6YFfXlCONF8WmBBcev
p/0Q+o7y60Y9aJwnZxtyLh6AMrWqvb5aHGUuvGnq4DqNs/ztkneB3grLj/53Jw7rWIjl6lrw8wtd
+eNam2Z7UZd+ElSVQwlVMIwAvqko43b1g+a0hI3+LUOzRtCoIhv7GyFCLhqW/0hSxdl5/EEJIYA4
syzzaiGycsklh6o85Y5uqL2Y5KPYBVWLckKk4hmRId718de4dhDPtK8RBwXE4u5DP8G/9PYsDEgn
JAYPXMFaoOg73AVsJGz37SZob0Cb8K4zkqdw7OlKn63rZhJgKvOAlZ+lB8p63Z482p73d/F6WYov
BrOpNlZntD35MERPhkESVEX/tj51AbvMWvP9Q/3168FPbeocFyytYdhgtVafth66pDnpB1ZywLgs
g1RnvdJegVw+kZdCJf19L+nYXnlGCDYWvIX73MZif9QI8Y3VZellNkrawjwquGZQDulLyeF9hoSo
mRnnMOmwz42rC2NkUhFFy/4sLVWJMgDsyhHZiR0DblEQcx4jaDNYiSTSx0/QoORlxdYxCPAfw9KL
zk2XUSxCDZDzBJy61HF1qjR7hyYxB4AET3Zl7u0cagucNUPflNaEycRZYqo+BUwAFgCK1XTm+Qv9
A0URKkENxG7oE7+2/njMo9n5Xd6afatgyYNX61v6EYQ5DhNZukTaL4pmv2UzrI062e2jO2GHtw6A
+svR8LK6kKiFZo6/7bu9cu2tIjvNt2oZdA8wRf1JUeTv+QGCm942bY92txLuUuziT2wDYUIoUCpa
rbVeowTHqaPSmOCe5npixx1SjEDCCYn1jnVKebFxZmLkQmDON8WlRti4m1DBJzMvNV4uo0wZ+pv1
w27YAzo8BOZPMwudHBuetzDbOT3tbjcJef1DP5m6pGRsiduFRBXkq11hgKU1BONJzI/13Ehn5IUu
NomMOYRp3mhkEYtA64U9ln4eD7ph4pHRADnXWoRVY7tO1yNETkKCHIRV8qzZ9wWFJW6+kT5rd1Ab
KEITOfH09L+w6DcRT9lBHOBiznj9GiXR1ZGG/2qwRnvRzbIxVUp9F8Lj9781ciLoS6T3WmKNDjdG
aX+2le69u50JJ7Qu/5ty/FVoKfScvoA6r5PrOGeMRY3m1BNUM7vSbUOF9yuuo4TmDPq3nY8acdvG
IWrVWCyfhRf8zHh0NybPMc4eBrl+Kf8RaDMmwxfWccETN9VL3DaBgMUJy71vipoQUW5Ln4SyVwsF
d/nb6WNEJD3B1V/eIc3CINf6wW3kF9I2o5mMnlYiWSd0KqvMfFS7fMgsczjAld2klc8tvJ10sh91
zWlhYg54r4uE8ChZ69az7Qe+rYwIImO4PiE1vYoqMmlqzd1rWcz7mNR/uqDSCQKn6/oKam7Fg8So
erLGBAG2MIAr2XfuTiUfOY3E2vIUWwe4gZ8inxstV0PpAGbRMKExu46jHI5jQ9dp02ryFAx1gkSD
zN+sIJtky4+IX0nGsyAuoVflTDywczjpKLmaDq8S2r3iV7AxhsTAUfP0FuX6dAeSVU1HDhFRmZlc
WU1hjluZUOf9LKIJ4OvbKTxUTPSnhnW/4hZW9KOJCAOdNgJH50QF8ZMyCH8JGGV8V7xG6Fp/fRrf
o1vAbIYK8d+IKdvGXexIv0Tv8BgqLPRnhg+6y7R7JseOZYefxyIGY/qBa8deq68e7old+uDehsXR
FwQct3+mD9OLnFKhuHMss2IQYumeJ4k8HfTHWE1foLtvw64TSrzmkTQUDLooIf3T/lMiflHznA4e
pwzkawX+EXtA7f1oYX8Y2xhYhssjGwhABmiVcumsxmqwGWes63Ey9BIiFrLDKqPVO2blqXNPSnjl
Zczye7BdO1992FYSb+svZypkmfFeOKkhY8OtIjkYYejhNKwl+XI/u8Q8Cyeq4OFxjhiEMfLrAo9n
YXBxkzp2czsNkukiTWnu14lBBcDSK6H7zeObOYW6hCpW8XRscTPQQXXS3NqBH4hf/o/2JecUJNxO
x+9vtl5k1d6EX0O9RRahO+zJZp+7Zyr8N0Ishj+lyj9oomhimvzIsN3CYNXlIBh57peSLs/ajOHU
eyf4GlXDFsVmGxw7gq9XvTRWB7RyjQtemI0CEwJ+Nb/qPcFUVKVPc47H8mt1lsuf6O4EmIfIG0x9
1oLiLlvnP7MDDwU213L4UPNt90i2MuhJSvrSgkLbNcJjYYQa2ItoJKY7xWYjtsmFal0wz/L1ZwIG
tw1VgRqOOVx07clU8rIm26eFtvDtwv1WMH3oD5Vzn6PYKGILXbTXwbEYO0fjaxhB5bqVcmM7Qj/1
3D5fqhD2WwUL/qcR9/agjyiZZfU2DyejhfBWtzVKEPZFjeJ8Es855oPqBxBq5kqADi7dUmObiyBU
h1Q9Db2Ghl2If8E3ATXhEEphmtLxGg7WasfHrPNJClENpxNra+Ubg0nHQq9uPjXd/Jp+n9xL+VcZ
lEHsjCloo68SOmzNHlmBgsYOEtBnJB2hARVLWrXRQxVfKRyKh3YQk1vIr0YUrrfUl8sBiy4/4K4P
4v4QwdiThd8+B3rUGGTWLsaSVwIiCYJFJ0UpnjB8NbP6sgMjVi2Z9LaI2UJuJbXssKYqdvjfUPL9
okXZAhe9KUF0orHHo7VDJzL+KUoY2xPzkT74VbwHmH04GwN195kvbFGhigmHB2i+7JK0kzOg7mDD
0btqILkbXPnPQVYTE1qc8Bp54nFkoN5x6w7JPIrkNStm0pULZYXqceJ00Lgq97WXklFtg4bSsMLC
f5Lk6P3/LMo8T9TMwbPmQTc+dd5lxF4i0+dqN0JyiFKZpeCBawSgFn46k3BXJT6Z8BezJwgIYbZ4
G0qfJOqPhGULS9KR6KRyKhWjvKQyyInNUqxCX13GRtyoRdnSkmfR2FQWkqLGLCBObUZYfrb7gGJt
/YVb5Y21xsLT9skswmV4fN5NYbrtcsfpf/eVH6YmOExTV4chNHUeUSPCAyYW4lc9Z9Rk4zYVlHMF
7GgbaPr8lUO+yVAwtvhxVbLzRks8jNHJvEfN3NZ02LtKrpBaOi8NQdwL6cVv7LiFESmno+zUN5I7
Qe52UeHCZwfzpF69ADcXQ1PItnWHL+DZejG9Kw2xTFdAuT2vKRdSMJ1YuxTd68uE7eUiWJPP4yII
RtRfJN1puz/anED+AtJ1DnGG3DaqGdbzOoGSwLEO6//hRl/zT4Pmaa5dqOucjrRfSzWBeNfI9YoU
uUGnDEXF6MhUFv8EcjeTfyYCJJ90c4xDHNjfEUK3GWotW0qCSLGV6DeZodUEo/1szf6cQP0nKN3T
ejChZpudntGUbtq/9RCWXI0Qa8WRQuiY5sHnl/gyZL7IA56g9xWI4sl/VjGwBaL3Varnx+UbnrCh
Z+pzJoIii8HHMVAI7oTv5S2NNcpanFKKcVUc9jHYJ/+NEPKY4Seb5cX7ApKqgbrbwkwbNhIhElbk
qVI4jZjgHC1rm6859zdOA+6fCQz9bZq1eSb89Wblwi2hTCnPGode/9clfzuEittcwZ4USaj5xdXk
yL9iZJP7VB/Nw/lWO7NG0psvD9SgZNIT8nAoD/CHD0c3vtQwACwjR0dLitff/lvDoiE1Jah35pCk
oA4EcJTsar4EjmoriftgGyf1vxA6b5XBT+us95HImLfParQ+EspOkLDMUNaJKsghAUzTkrpPzmDg
evTETLdh/eFSsnaNthyjmZHL/vsVpdqBK/C/miTlMBfuyPPwDbXhgCOJZrV6wd9VwCDo9dsiF46w
xTaAGuoJf2Q5QPlB+T/Yiw24LPIwwd11rFraHvRgwvEhItsAdwv0iPVGYgVpJXjyPEHWKJsSgcSn
qziD8TevPinWzjfzKjdAZilmjgS08u4kI0OUZfsND3hz+TlJL8QMFatsR9d3fFdxm6JB9+W9+BE+
E1bCkpH1tZMhQ5BooP8MJ+o0rI7qe/p3nJ++ftBQ4WvedSZLmFCJm7O8frqquvrrebewzBdzeIee
OZWjetONvfsm6xPqkVJCmVXBsRLDrsD1PmEvJtnA+63njnXv2bZeAJHwWNkos5NFAhRe7AuDRJvt
QEtuFi+P5AwINGV6iWlmi4Wr/bu49MHbsQfv8K60YMzdSH6J3h9Ed23W3MWlVKTn+L7l6kE/CU+e
A2Y4Y9y8KuNZGkLB1oloG3rhkxTZskhxghITbx1GjeQLLE4gE6i7NI9Ikb3+zj/XWybNaK5MeEtK
hBECXl/dLuLeggQBZwAY4YNO7ND26FXWyxf5BiVX/DZjKOpRdIjRemu2MWbKGrL/+Z2ZkVNf31OE
Zc5iILfvv6aixLbbLi4FzZiyqkg3HwURkiTrphgMM5z17pobZynD+UBenLyk2h2/yS3E3S0pJs9R
H4S01umO5SXmRlWxYr9YabVH9ButGkjHj8JaJ0OiR/n4LTb9mlYOhJBNMqVI3Ivocq11tuYUf8nt
Z99xF9YSER29bt4+z0Lwr8ytt3cpmfkD2hx9l98k/zvDSD+r7x/z+WHJShPmwRDc/W/Djdjz+wMH
NxQEuAKwOI0uA1wcry76X5/PYrCq6z11QkTRVj+aFE8tl1/hl/8w5zEWhnTOIbItvjcpHLAb2B7b
qzoK4+o29ViwU9VKUraLX6I+J2QPgTccMEcxDlS10sja869H0vHI3yseOUF6zR5jKRU+kKnS2YZF
Sl3r0kbOJO3BqPWOse49SWnuesLqo8boBssh+7EC36ghgbPP8qvqCv6wZBspILujScKSuRFp1fJ5
7DrpKltit0Eqr4/7hy5aRdjg0mpXNyk9H3Lf0WO/NAFtblsFss3MvOB9uQu0LtpEITBSjc2zDl5C
dVdbMVpBpMwltbOkH+xXq4Yq/06HiZzJa0el9AdEsSG+xuvUW17K+VsJOCXvAFB+VwaGzEmBRGom
S6SNcT+3mvEpRgdWSK4ELGtX/06OCxc2difJPcfuSYVlmBUS17auuBweEb1NqK4xngwOj1YonxwI
kB6hSuoYLZV8Xs+Ta2+Tonjr/WZZpvFaDOvt2OlwweGU0AMgHauwKdZbW+FtJYibqJfaNhc4/pMP
8/ph3ks/iKiCJ2TyS0De7HupkYtwE30Ady1zsDvraojWA4vH7zNXsgZo+IFK6UH+lrnOCt2nLyMG
59iWIhgvnMI/cY1dfaMMBFr5uF4OQyUua8IQEbkFp1oEC5Rvcis0FxGXsqyGeUIuBhqsIum4Wgsv
nE8g6kZ+ndTF3DYbeLXxE2kElN8fxFk5TWiDEpKaLQ1mJbF94UtcOQXDWljaiYPstnP79YChUceW
pJlP0b2JTO8JtkAqzX6XszbABz/57cHd/b9qUuXQKwpumkqCEhlJMZ1B+iuiZe4FLZ9uniuEqc9u
PS/9X5yb798yUfNlWdDxfYL4JTXVLCjLD9IK+PtBOYYNSFs6vTvmaFgCYINBNKCyhbZs5XRqRvEK
kLinYi5DEEmAAIf2PgGOtG8iOJbnSXxfIbbZRCZY6UWeXB6CqOczRB2V05GU9rxFdjfIec33SpLR
sxe1xwwK1jXVPOoeH9DVmx3McWB5Fn6JNjNuqZtd7Jf97mYAsjuaDKovtj62L2dY9cknoF4uT1m3
QsLUGaqSGW5sToX461p+y0HziUhwojq8yCDG9J59XT/PdpNzJRRHXs7JPryOvpCfuv0YINClnLuT
AfDxfWDOc+cUpLnm994pIpSffPDXKqovF2g/e8YKyGb2jwJ2WFp/kly+2L861+CXNl3K163kBnQB
2kiUTVzB2+ySpS2kAqAObE7phYDyZyfeUFpqyyUL/gvHNDPfBz336Ne18SzXKWQ9BiV3r70Cv7I9
wfsAqazWV5jG6qIZyn1G/jEVl97MIott1HYn7hNj3U3FFbpSob8jAjJMeeXmgOqps1HUdks3ygFI
C0pyXghuB2B9oZ+q+8bnqHfcd/eBvuQjkynkyxX3nRVuoFN4i5nMDQno5wCea5kCmkDD8WF68nus
bTGHDxmq3a0pw22iPxQT/b3SDBucMiUvIYx/VkwB0slyLPT+8uDBmu+gtUM7nG4ER26EQVK4NdTZ
oAme4eVZ1hjZMRXgC8OYxvj/D9x+TmmBbjH3cT0xjfTjzmj4tq+WXwU+UBChcekhmt4k68yU2DcH
IOJn302/jx3BmibjmH/zyTSAgMAzqnrJ3zcCDGfpbQYQ1cXScaxNJT9mWj30MdFrX3V1mGagYUlw
zPLMNzHpopb2/MG4bdLDpb4IjERBg5bW4TSyd9T5B4EMFqnzKylWGK/hwkeHbOQthcjaelfVWBvu
dxX4OYAatDaeVs+Qp1Eb+DdvXwfbcsYR/KL9eutSIqtzSRk0NTchY4nM1oiaTHl8ydZPXkx0xZ5q
5wQtphG5r4blLjg1RDK3XtOUuO8Dg9JKeC5DqqiUiW2dLfOwQ6forXLeqMGknaE0Jrs1Z+sbleh0
PCUJty4ALCwwUjlVGgm8R1RAUaNfocs61Wktf4lB36oM56Jkq0RQOZFrd2VISqxNJ6Dnmsl59AYx
pTxJPDYf7vA8qo5o/eTIOWp/LIsSamAgfIf/29Vl9DR2SmapQZ0N2Waj2xLASvzenIkk5OijcAKw
xSAKBaqlG+RRbgmcbxKtB0H5t+ETsrsUkwsa4cikAxreHSi/KKmrzEOr75a8kfspf2IBKNUgkPee
PzG9RMSWpVbCtR5ow/Y1BlnD8/kBPwgoLOj5+i4HLysC2vLSRnbPB1CaNSgdaai9pPlbiWWY2m2n
vMOSytjVLSV463+FXodlZsBU5P2zak8Si+6mQXZufqB/IlQgP63i1l+WbwS5K3rKMEEInI44fFSJ
SCPlBc+G2wqWjOrfoVBhrutEwYz02q6as0phmiVwOYzMGmm9DyfyhLGi+XxWIMxnQ8/+mS77POzH
csHw7iNXDqY1xU+bFpxqWotiURhE96mJDTrzQLREboAJSPI5TVZnMV6P+gkVZ1yuPgqzX4H3Mu1j
6Q4FaSngxpApSEfsm6mp86ISZ+PbDuL17vplki9f7qqiQ8K1lXcchhCAIhMPgPUa+JZJXUn+vS6s
556OeMiSrxtQW1sFI/S1GETo6vjPdOYNtqmuBV7yLeZLzKZj+jee+TuEVoFX7ZZdCCfY+CqGUxqz
zMItmOlAPwNuYNr9iOQKzQbE/qJr7rknfB77UbfRW3Po+TRd+87s6ssPLOULUWGzdJSyPl0FK5Kk
W2Zl7JjvOfu9Ad8e0SNgWhsD0wHmS6LGqmrxf7Kwr+1bftMrwC02cufsXYSqUciyOEix9RHK4xTt
GyvqgwKN1hJQTnsb2VoBaBZYybvLDRb6bB8aztslN6u7B6BsgYG5iduseR5BnOnThxGdBDaJZnt2
45NvX+fsZaiDRFRd2QSAS8f7tRusLMZFyt1RhLs7gGw0Uz8w+bCW/91vnPefjb0ENen3yZEhiaV9
MN1Hbsed2zbHVZK/d6iLVCmc7j81oakCBUbNUD9UgbtyWIhV2OvUmXwDHGzg88Tuq20a5XcYUz+w
ux4BYSdg/GTRKY8EiLqRR2ZH8pjbRDdfsKLGZMRevVKIa2KskBnaUrgXUOm+zqY4WrU8ok30giDV
a17hESeYZpdB1cIgWJkP7kgF8KxybREPGmyGh6LiWdtNWWho55yTNOf5nWNaU8TqG/bMQfBj4zH/
gB3nE+Do9oSM8jfBXmG54daOnEKEEQVpRu05b/KDWXZbXw2s4Lt1dPAp+L6QZfE5RT1zh/PMq3d2
iRGThT1Yto6GfGiiNH7GPZB7OBbsQ1Tl6QnIQ2dLfhOVjmPI32Rc4QW2ccLsu9DQhh/6gDYY+BJw
cvwpYRi5lEIX+7vYewYSn+gG6IeQiFor6dXWhLLVr3wb78uWA1SbEIU5JMqq9DQhPxODUW6sZjaE
Qh8rA6ans1tEbDbL0b4qXgw7lM226zBzjP54vjJzUHx/qc1GjAUo5kzMYmR+bX9ekmuvOyA0jjQ5
fTtAUIGSPLcRhNXPxLe7ZNnxST4O0XG1ZU2rgoXk3xPz/Hl4VhLjjxSrmRxcgSaEusa1PKUEOVwV
Z08DomoCcF1OmXXUAXr6l4AAcaoc+jAkjYq9otJoogosiGC+rd3RLZfmEpCgSJX/kqAw9QGV3OLk
4ckAnRdsHdMURt3YKbetl2ByRXB43pybcCtldaOQOMm3YaEQoifRmSw57PH1oUtR6BdY1hSwr1lu
7A7PHRfcKwX+jYJ+MvmgjkRr9d+2/77Nc1n7ORVk9680DFIAhNr8IliokCnsSSb9LZnCJxG+tOa1
FKp0HYVQv4TKcG+zfZgMsZjT6bAy5W89AD1KeQ+/63DsYvfdnkqIgaSTU/YE/x7WyKeKczNwh9Bl
qogYjcJvA2ZgC0JdViqTpDC6yhM89NNyZDc1urRU3ofOy+yIRJZr9RKLCcwWxnB+ecdslW1Nk0tA
z9sso9b6Ak0pJFChFLmvx5KzbizHMuwI9oOZJB/RbWhuQuO0mSUvEdWoK2CcP1s70z6OQ6PIAA2p
HObG3vsSfOvceElnvNvbr6QHDEy4kq0yB2DjWpCMajIR4THtBjnsV0Kpym9zIxk6+BwTqWIeBVHq
5UdSiPzz/e3YbIjXecyU4/Oyl8ZrpSMUYHMHVVCdxoap3uMoHXbYdbFyC5j6wvO4wVadFeNQnwzA
A2q4yaiBiIcTzgeTxYCa0DCAQ7gNChT8vhocPagrYW7pPj27q4gPb3d+/H+XjWIqgF3ZiLdtCdgP
fPxVNsIiMnr7XJJIILTP7KJmcDZWSlYepf2H/1+ks5zI2hmQK3cAG60ji0Hgzw1D3LrlHnJxZRQ3
tM7bM4vLHnNu+QkTbbcewpa2QYV0Hy0Y2fPTP+MF9L3hcB2kZkwYwYwMCGy9Chj9omsRsWnx3tNH
d7rWTBE1jG4yt6iT52oESgErNS9VlXtDhQE+5dSfC6LzDRg6deTm+z3ByUR/P35rg9dfX75q/R1C
A/IZb45YpBd7+mliDM1POko+og3OBoFhKWCLqsVvGLpDd3LROFg7LI5jSHQi9NEYlAAVk+/lgzBu
bi8hCUny67UfMI8GBYb90IBAR9UyyIw0JITHbe/J6EJfiQ2NqHdkywiyiuVZ+VBzQM0SG/rvRlWL
puMiHpAdzWYhJMr1nRqgjDOStliIcV0PkooqWL+IP0s7gZnYWsGt0E00kwHlWy5FMrPzyzO7THnR
GDhBzxSfg2CyFhEgEDdjm75dbvnzg3hlbQRD7F2was9WIhPDxYjEkl/eSbRCX+dAEVIgxCFd6aMQ
v60crHFgCh1QrgNRkNNwieEAGocqDCq+cot79ENxP5BQx5JRvuVr+q0qd+ra/QRBwfBap4Kab9yS
v81BVIUGQ0L3yzArkSUHceGolHlL35WmobNjzQyWgJ/zM2aWSBU/c56gSfzdrqvu24FAPc4bOS9W
0IEbPqkYi6WTMJqHJUwbkeNPPT7ez148vCx0djGUJjxcNTmJWV0dCS4yr2lkwwKMjzwQC+gBIrjd
KLHO9pC6wcqpCqOZLWTPT/MRHK8QzRdZT2Qqnt8vsDpw23hFfO6XCEqmCNz6ZjNAZbulu3pPjhXG
lWNg7Wu6+PW4LZKzNLMOAkMDescPSsOGyCcj9JLXjx1/AvHLbcXSKtrO33J0agiSTemGD/lCotYu
IKtDaGs5MN4Cw1FIkHdFWtTRaFEom6GFW2YjjahDqJ8bEjydKQDB5IJV5J1ZszMUgsy2andRbrPc
aQ/u7k0FY6+EI2s9h9rBz8aZYb01g3rRNoQAkvZxXZWkvZWkN5iqOWMMHDsPmsuI0QdLTK/c6jT8
i+oE0HZSiEPJYoHD65yYa0aK9ySvQwpdhQb8fLH0vDf+LsQ0lIIQ9HywCZRamlx5pwPuyuvSpOQO
yi5ICZo11Cf/q89IKrSeeXD6NcprjippELWHTwLuZl9V3BByRubbZyLx0eplFHkBQPfxs+Lsc2vw
GR1AVWTv9sjsJtez0gIvp7tNa8J/ngXb2/QEWJx0NNqtWbR/fdchTgKH2l/UNj556JUkR2vSYdCQ
0+Us6M1xYsF2v82dDShduFgucc6OYUig60CB/dI+vp+Z10DxTVs0VL4gcPqZECApYVEXP43YNbPU
6Tz1/aeeDvf6G2AKysQw8wjZ4wwuvd2MRs9RZX8b1vWNRS2C9OMF1bXPXNw1KvJ+wVcmRiE7aP2c
yMKJqIDgx3tJ7Lw9jmlm210RxHs1LWOpl73eOX+E+X1FfuXnjJHJteNtTNhHhdG8VADPt+JynQMk
nsyW9wmz+YZcc2K2WVGEeDv8iUXRGnOmKW+8K9A83gMRe7PRTJOqcXw+KTMq1nyn9G9O7Yo+hidY
iduwtk+Zn/pMUnngWnDaZu8rxbXldJPqZ+MPEDg6rupykpaxYSfsaYdpBaANf/bjVB3Ox/BQfYHO
a95SQFHpyBFsDazHQ4+onKx3GDGJe25kPYPGrHJzSlphMZk8CExc8DoAV+nFCrNugh0M5szOdAdv
1sYrcfs1V7S4ajP1shCNp7Vi6STC0lcKUgaRZvh2+vG5w05+wwZD+rxBf/PU3Ci+rW266gRXk1ep
/SVKooltobida8HwrwN+wQvJdFmOggGzv5jwgdTKGgkCoJh34yR+zmSEb8C4isiv+tITU7E+AvVr
SLAatTypK4ulPj6+B2HinPgN4fWbP9fXQ//mINXNiLvwqt40fpNIJ6EMoJ+3CALYSHjOiHPEWCWY
ueJW3u1uMuu/kYsJT4e9j9ehvXezvoRwhyuC60HekSl6nKtemkpUsQ85sAR1BoifpbXqE1X3/vkI
PaAukXdlP4552MKaZz93GLZkA5bKqeLIPXJUb/+DEvLBTNnM1bsLA5MT1ptyCXEkmu5a+2Dx15en
ivEIZaH8veSKaUD7R/qR8xEh7gzO9C0xc0zQqqZyQqbuA3UPVN87UXVZsZCavNWJCiGhEXim54fV
188V6VaNEsXgIhH3VazMUuDFSFB9BQuzYCp5Rhn9ioMXlK9me6SA+3WhT8xbtYED5b/HBpQGRW6p
4q5EI6X7ev+sON54viSTxHIJvKZ5h76Du2dnlr2Th2neRJFMpPQrICizt5LbVrN24gXqh0bO6kjS
3nZun3hQ0ytj2B/D1skRE1ddW3P8z3I5FvYzmuR4+erwhG8hSJIeYNjNtyq7FHxlrrZnlevmJccG
A/sZgP4MmA+dflFLSY0zRrPAPsKBhV7/h4ooK62Vqx2Bt/ZrI5fpEdaDgSXsxHGIb1pN2PeT3eGK
noUgCfrLtQaRvfvYqTUvpnfjynRDTO9SXdllhyOIbYdisvMsmP6jaErhyH8H0iEj567O0r94BHB1
mHCVLtF7y4pRfG3fR96i4ce4yEMTY9nYjJhRqN2hTK3NoKHAnhUJ0YrfdRebJzq7I+tQhGfhIED8
qkgnSY5jLaGMccmob+48oi8FiTeWz1SF3ZzU7umHWAWfq6JEnBfY56Giq7kc0koZkBHzslg3lNA4
ooLF00PE5fiNu4ru/SQyMPjXKwhglyKQaCy7xlzQTwi75RGS+quzPDH/d3tkz1Fl+wxlz/BI5tW7
RtqczG2KSXSLOBNyFj33bnC//1zihxp7k13iHxccznS/qtoLDkmR9GshZ12BkW29CQIldgSa7Dxr
sNNXFFVAJHCTj2uHigUa/Q4pu4LRYKT+Y9+Cmhx9/IfB0yOKBn07yHX14blysgft8baDFo/JIsHJ
hWUvdlsrEz63UqzTw0DESVxVWC/B6dkrdz//+6WlALsvE1HGDlBg3MqAuFHBcTfQRyQnxYuYlMPl
tAJhhHClSlsQ8p68cy7A9ZuvXWfI2A9UyJ3SJjxrYQq8Zl+fApAZCfbN38qgxZ2QM3iAwly2StoF
ado5nCSQfasn8cMnm64Pt90nVFRlnZlv/j/H4qTu1kia6JyqPB0GSIsWvAqXV8C+3UzAf0oba/qT
4zdK9xHz/ZT1jZ7YQmabIeCe8lm3hO3dN6YfoUT1nISPWSjW9ugG2Sqa5wzIkL4SXNVvTUKKomcr
AW7KNlc9hdVc8NR9nqS9rRzqTen6zAcFTVYzMVSS3yK2tY0kIkcav2sx9PEqHUcVftBw9YIWMDST
dkri4GcqHtS6Pwunu8wFdeDAxEp/0r4M5KSINYBEpSH1SMPu5A0IUQvc8p7hrozP8KfL1nZbTSmQ
okuYMRiS/pC0snlq9hZn4Rd2x7sjLbawroAlNVNEEvxNTPVevmjXSwveINfYXtrFOaeWdWhZIX87
CoKw6slroQmAPDZcZlXCrW1y/R/49Y/FRi40cwi0fty9rYRs++cltbYyuZ/ZcVUNT8/JSB9O5YFm
wi5rQir86c877LsiVHR9GUzmOy+tYAhutiNHEzKQzjC0S1c+2jWJbsFmjiDu7WNekB+AnDUvXkpm
qd9cTOenifmavGDqf/qSMDhZYg3UHxy9ZXzCvaZSa/wnmTTfli5cftDnYE6mk62TZcpodjlRT6QG
9OrqFZ5UW+g9wD2EA4xcZcgmofvepivy9U7X0MXwS4yRmzrs62YdxKxZPKuuPwW9+mQQ1Ckke4RC
d9mAQGyl+0Srvvg1b0qCbdkgi9l+29UP/Ki92Pr0O1B4nhW8VVb30a26XxqVETGsTxjTZersUNcM
XAYeJjT8cYrwJqzp9FJRCEOKPL3BDQ3McCauZAvjbVdAWKS1aKehAkTVk9VCIJXbM2ofVH9SprI1
/xy298/CBQpZsX7Vpa+Jvo9sUAqqrDrBQIl5fls1sJml9kgcHI+aZB24WYtvxtJP1iHpZmfN19Tw
NfkzRyIiBDaRXDIh0QrPFwtVfaVQsSeBQXE7YH3CaVu7vNSkz/CvOL+5B9ZPiNrcYlNRpuTwEvog
MQlu+y8KzO6gYikLFdN+TnYBXIxFx3IP+p4vr7sFkYxaCk7M1CPfLRroXlQQ3b7YusnXnD5Y2alN
ykWgTyDHkcpPTlSrnSb5gAR7Yp/2EUa3Ln+D23FHlPNSSzTLoZzd+QK+v2zJ6JxLWGIu/urbs4ke
HO3TN3sSuR7MSi8gNwGDHhxXJ1E0gD1YKhgy8gH3d9tlM+uA/eGlmnI505obNph5+lBY+YVi6Nth
eDX0s02Pz20/uPw1c8nyo0YfHcj7xSVOW39mqnjXkyzWrHq54DK8NTwi9oZ7yu8nvjiIbC26TUE+
fOdWt8RE7DjqG9sK73lbu7fk8Cnu+bGemO8am12BZsToM1NFpSDld5tVSJrpil5tilI1WchYq7z6
IMAYCBp6lb8j3khoxS8h0CmuWiu35E+tmGElHZ1//DHJ2o8aHwrUz6X4UjXIgYScGOC+ABPDwHyi
zvcRabkO63ikIOEa1+HuIOcONouVuy2i7nzyi4zPXnlMIfFgmIt9vSyNMClwFRsfp3VPGvQmOgyx
F613QidedADV7MBG4LPBAa5SWStb54S2bEp6I5N0JfzDthb601SlgRRx7Hnz05LLeATjEMDT6/Gs
vkDUigNyDhJ5hfV9mjVe979I0dqmAMke5f4LYDiTIUN7iYJAOI+cgbjaLGDnAaVsHcypmtKJbxkF
okAVQA2SbLqaAEamDTe4mYOsqy30I9E1ybm8i7i+b2uleD9tbJzbkMRYpgJOT5WzW7azxT+CXxQy
DYFONYCMpnOD/Mu9omceDvvKpm6baXEjaR1WxVfkeOwUK8XNHiTM0c/2jthJf6lh8p5B6qBe8xfX
Hb4Hbiyj4tEp2bhMNS0/h4LBcQSJzikkp4ppdmoepN9l9KhPyhla/oThwKZnjvOjscnq/oHa3N/K
peVuZPT1UbIE84vvoBqV9Iv3k/ToFEiJ60Bokhf3Ebm6Z6/guIjKCYNM1DKphhSf3UjdYY9b4SB7
jG6u6R2reoqIaSVq/ae7gDs12XroX17YEnWxEynR+1rUCS59gOw4sJVz1BHPnNuw9VBDGNSG0qNp
bIXZ7P7atPLWXJv7y6HXnSY6AgmME3b1z6Fju6oMZEa+EcNac7YQbb/uka3Y6IqaHmBG3ILCRJj1
YUEqLZNpomXzDctBBkFXP56tMa5Y1wpUKdxQBaZEH48S530Iu2XWt7xVvHpgG1fthJiNUc28AMbH
1OK4A1S7lpxbxDLt3suvPKbWVr8BRQ5x+rZTYDD70vzQZcvAIup1d6cxhgDvRT3llq4VY+Oevgg6
W3F6B3jhsWkFXedR0AJlwyP8KAN+bHwJ1JquL2dvWpfSH0c8HoXUxJCvO7tpxn4y+2KNTRMwK3/L
HpCmBTKTPiOm7nzCxy5fjmkMQ+mA8Ed3SOp9L8tVTDeJ26P/CXn430d28l0ZOKUldtAL23itak+K
CRBL0IAYLWP8NpwH2eDkyZWUouGVKuLG4y+p7vDsyE9rj+s89E4HVUYD7RXw84KxZBHYDPME5Mne
5Vx3g0Yy7RUwAM9ugX6aqPIdnV405tvg5zYwlgft8XL2ccmvrx0ew00aEs+bP2TSIQjRuQLhXv0K
9CkGVJDwTWRvyjfSETrgKA3Xwi8k93cuUtbhOX4K4N3S3MDElykDudrHfzibHZB7sXgYyuyP1QMr
cGKKlcijm+JoZEo5zqPOZWHduo9wGi2z5JbwivOnSXTketliZlKFk9nWnh31DJnTsTsrhA/BjcaG
Zcs6Ekt0loBEx0JNpvcTWdQzXW6ELg4sU0Syqh2T+eEJYTam65Ov+5T7E/bsoEnyoqIP/3hXaeSM
Nz7I4bCrwi+h33GSAZGCNrDXsOJFOlbFQRuAX07hrAPI/vKkozsMUVmsWxbKwJdO78B0pZHS0Ibs
An9VPK63NmHN574rcWvFIfAKl2tP5e8yUlVWian1Iaqwh4I8qx2pwqf+kzim9GQI89vmly3qYURo
NsOkIqMY94weKSS7pWfUPgz34DnpvqRvpbhCx8GUCiiYN/mi8mwsfeM1cKfObuHcMRnCv8Wc0WEl
uKfQk+BYnlssmv7l4FGYt3Z1sy2GtHgSvkCsTCuLfJqGrV/khpq8SoxgGyc8QCHuI6d3OG4OlPuh
qNIPgsHQ544h5teZADcJbtoHxw/jU9clpQdH0copjHOmM3hArYeNg6ipLfyMBIUBLShgKEUJEOIz
LK7ypPPjPh0AEHXEVLKOOHzTTL5CMPTsXP0Q54S4ZiGo8jHyolZlGjNltrygI7cT0GNArNhVtVYw
VltxuqsWM9KbAQY81pWYuY2zG87mW0NyLJTYSlXe0LeZg3XJnH3aFWAl9cuWkIohj7LkFbPgo8wQ
U+Wc7XtFpYydbiksQRxvYI3bawK+t32PfYgXXDiZLg+BwuWin5ZAi0UNHAXL2V4+izWv30Xvhi9U
rad9699Qk5bClGnfF4a9Z88Dxppv+w5NEVX9V3nNpg/52/6qIPvHpmrjfphSHpDIt5ixbMRZFi7F
1G8kli6ocpTcayUOEQbq0w7/85XdqdCxBA/GGXvpWgwow1Mcri+VE+bkSCPnYDeccAJVldq9amee
3c0jPTFadHZ+do+rI1flb0sL5l7E/t/X+D8HTmQoasHQnWqniWx2V/sS9WqZFXTwlvTIr9bLREV2
DG3jg27DYU9rmksGbqm1sNQIdR2dKdaLsaUFE07Ei2fOoYQvfPdCVDRpJs/R26ANDeoAVOY04+bH
ZAJo5LSKOL3oPDk9HQCxnRMTDh7QquYC3YHQalSVdGF0o2S4ePQx/j84inLNSodjnqMrORnL2cZt
rDIzWDwXrtk616PxtoNOrJ8nzzRgW5TfbGhHp6GloMu1rWpgXMWgN32l6dFodYtk+ycU/4yTobF1
7opv62uoJRPa/uOBCRFmYkqOg99alXs+JchloPtPkTmYcB206DaBUpgcKFzOGen7omUKp1AazIa7
j++KB6urXJ4SI/rLvBnr0tLbx2iPMHLHTlUbUs7uP68C2YIoeIM+rpgIk1UOCOm0JKikDumpw1oc
RgPZWhp935NCQckHSCTJtI3s8fo3HbRfyqyamFXj+feE1Sn4lrt0WEt9iPAxAml/fa9bgBhkWhG7
0sVz1DYbfRe3nQZtC+ns2Wke8Bflfd2Q/+pC6NblETDvLiKPAggfBxpxAfDXYR8AnHWICe6cvjS9
Ari/h+RtaQXEn22cwjHi+9hn0aciL4VAA7Msy+3cq6NKmAxeEukOCM85W/Nrv8t7YXB6mmp7dQm5
fmp1+DauqxgnMYGAqfLTeIyLRP9BpMPYgm065qvmAkT/1tSAbuuluxuU32HDZmZucUosQMYvE8qx
k3mwy2S0PQiep0hY6d5omq3seI0dhedk09aNwhYbb1Z68TFUu07Eahs/6J5KMwdZUl1HPA9T/DxA
UzJluzcs08+vRNEBdvKETsBnnkZsKNhqxIhqhuFNrSJN31V9K64Qe0mwTvBqWbALOVb7MT+k1L29
cS6uHHRBMl4gWE9FQPMB15SQMNBK08EEw8HYYq33wOOUdMDQpIaYDwW0CuP1rssU0rVT6lOAXOQp
ZP0jdHBMHVpawQPMp1/8O1HxZVZ8NoM7NXp5HD+IxqLB4I+XLdZJDUeyReIwlauxXctp5jJGMpcU
MMIdKmmddBKv2hfAd5WlS/2qPAo9n199c5RGiWLHjTY8MXkrBkmm8j/+Znp/c3zwlZWfQaQDAeY7
DJtfCrPCO5d23lga9r9Iq8U8+WLpNWr8vyxcoifctV3+8zmj/k/edcREe7EKOmdaHE5SGRhsuj9z
O7WxgX9GHYRUQzD2fmG0ui+M6rVn4w54hAoAnEWUG6ya0/UvnnEaYYmyevQRq8s3Jsr8lK3f0V9n
9MP7BIyi8/V9Y3U5/bIIGchFLUpordS6fnTyKZf6NX2FSXmwOnO4Mq2lB53rBpIo/TUtbivi6bCZ
mUjIS4Vb5lnoraUpK1hxJ9IecWkWTcSx8Z+A9wxu9Rt3MggzVk+UvpwI8V5nuxfdHAYQMz8CBF3J
kf8lpW7S5bzU0TWK44DD9KguRtbX5oxUFL3eVN+MV1uRG6EePp9JLqzcQ6JH9yBYp8gLdTy8pHix
JKKzbstRobj/xTZG0filGO9pN1nNDrvHFOFG0LjyZ9dEM4wRwm0UXUP6PIow5PjDyGjgzQMyGfwM
3NfOR/+Qx79ltYIJx+8WQvA+gR7DBUc1Pxupusx19JgTSxJ6M5aWSxckWWHfPSvTaYvb3Rjg7Hts
kzlNrJnCoGRAsfZKi91WbYO62l5Vtrg4ZRjPQk07ivBipI84IjQm9SU2juE++GZFjTFTtWJpgXyN
35DANzPQ3iXCEJUsfymb7kby+AykgKq2pa2kBK4HXGmEMWXyDrmEdoZs0/OKRIlg1sI0KxY5POA9
CkdcJwfOTFGwqo197utEhUsHEnA77vL3392FDeK69hMlyrp6fdYvgriTK/1efw85+w2JCwbEdpg5
sa6YWarWvA0VkndAEgCwaj8nMOWNWLLffYsEJHrh3fpGmLtAAb0GN1ruGDIxZO9wdYYpUBjxySPv
EdY+qO5qecgq0eLfdrvK9kSR4jwMPCGzDplP9xK4DI6l/xAM8T+amaZ5GNZ4GiL9F2LsBu7yNd2F
DB4Ez5RgIL68VuvhIcRAwBiSJxZu6DN1rZFcK26KHJnY6F63/9EeKZiO6Lber4qKyF3cZhC8eZIQ
KqRSXjNquA8GDctCspopp00IAhq56vTFdLhgrAS5k6yGMjPi2fv38BZJ2ovpa+pzLCskA+LFQENk
heHKivdlEprUrXqRkindQqByurPmEtuOkc7z9qnJRB3p+6aixsRqJPUmOFsKT59ZbI6CwTruuC3N
sCZamRaUBlO66rf5koFEYknVL605Ld7gWFK1rYBdBnk9bT/zaiHP4YN99OZVcpYyxK3DH+s/RFM9
zMr3TZPgaTReF0en8OeOGLVBm/ukyEQ309aRFaCEaBKCFeD+zPi3p9TURKFSPSUsd5y1eV0rpKvC
TB/TpK4MAtt//Z4ONicbnP8GUSo3jheMYMdE7BwuChqHhAOYnptRxpAvkOY8H1GyZfeW/1Ac7unf
GK24AaBZjnddyeh/rk8+pChPChWPSrNCVnYpDp+2SsmK6aFL7zk43vSPyQUiHNfJdNRwQ9dkARiy
be67x4JGcfH2GBitN9W71y4xDJ+6y/yUYb2Eu5BGoc7b5IA9VyMaM2WxvFDTD+m898dn4snUMHBf
4m51Fb5M8oLY0aY/aqr7a9oHRRfW1rowhwdHN+bQTWUf5AIitrgp2O/VXyraHPDLC1cYK0wDKnFO
btGa0ZxL0SIGHlaCU9ptaoq5F+cxjlP04SAnT1UY5bFmAsPQUKNHWkXtO/26n9nVW33xpYtO+FKM
RlcUFqzktkR2WD1XfkXROayXN8CbiCoWDTSI3RcH1AZYKEi39FE3kfvhhtwYgTua0ngR1+hbozl3
zFlP3/nxHPTtP+kGJF0n/YSQU+X+kTmoCJWVpuIPl69dLFpZsjiKDhm+v8C4X1VfKoosH3e3tkdo
8oV2esTFfguZRoqqr4t+6d4FPgjezJbltzZ8PQzuGbSyvRRHWskZGAnlDrI7hGeRRlA6+/+ZW+0Z
dMlbNR9alI680lFSl8hgzOn3aTTxctJzL5TAXrVzvqJz+W1+zpp1kHkEOhR2SownRWejWSdqHE1I
y4yulfchF1duvFrROuJqLFxjn1xZnQmhYcP5t5w6PnVEM/CmUYzE7jmVMdm3jJE3E7HPuYDzwZHw
OrLBOZx4XYabVi53teBD9ibyxi6fQlnJIF9iXhcFbYCD/j5beAl2LJorO/qMr1XZuqsyr8vj+Jrj
pC0+RVu7XGvh+O8iLrcAwE6JheSZBW8veJ8tyr6ofnVUSrbsbEvsUZ/2iw2zAza9wPr0GYpF7lIf
bIzoiXfrFxW8PIgPu1hUSo5Dt9h3wZU3uFr1P5CPUorks7xk78ZokxIS9RTuzr4qIaGXPIWk/M1d
6rBZqSyK4eCj/tvCqMVJSPGOuJqn4PtAfRYjSsiErOPhFIkBNwcvHdsG0DD0TY85x2GCtV0GAZ3I
OyT4+0ZMW3ZVEpwqiwfYkfBdxiT8EzExxyReZppJyItyH2UssdNYTQf1rYvm8841PJeLQQ3OfcQE
x3j1jB8E7rGjgDk2KpCf8nx6skIB1OS2ndXzTYto/HQ02yl+LwDJPcvk/r7Gh6YZBfr2C52xa5+P
xEeutXZRH49KVDNT0Ms0c/p3c4KkqZ1tsdeQesXt2JpGKMI4z7Y7+JkoQ7vYKqWx7+tLWnv6QL8q
qgjakNGPd2eSCp79zYcy2EVTW9KbZVm1ugfkiwCnWKtfvUYv75E7kP2pCbV+kiCK0QhuQV/y8mvm
Hcx0/F7RHXm/7I+R1njUwPIMydXiRwrlkc+cdZO2JrjD53mZhEKormSv0JDbdV3oQ4b6784PGMy9
9yhwjG6LPH8SfqdCpvGjO+Gwztn8vaGHWfShZ8uVFQiMfRaRGfQbqTChx7J9YMEPR+eg/JZEga0/
4P3ytUh3Gw527FkGEoJTlxFNXnrrCVvER0gxSB7M5J0gv7y46UUYfov6cbf02/S/Bi5841RcRHXk
OOvbIsHCkCXNdkGTc2zX4KGnLgD1fQK4R39//YwoBpiVWwTT2YuPzzLTPUwwAVVKugKb7bXUcJvB
ffIwgA+O/XGWSOagt/4CqGzftrtfqRE/esT1CBIALDqE0cSKGx5xwxiWwX0NY4nY3qz9sW+hSOxR
MFlJiXWh71noX1hx2eJZFRnc/YBl4oeuhHKZmcrtlzYq3rp7a2q1Zy+InvOYyFZ9wINo5YDgUaUZ
8yQQXhwUgIIUd935pUy0Yu+CdhxA8oiWguCvSixeqCS1pcfCiSfdD7dNWveuPrIUO2BpOO8i0Vh4
0nN27NhVEx9lcI/cBGsE6a6zf7t6L21zFvdHav+MZFF5mckM9KXKrD/DwgkOZff1WoC/UMqWLBUw
rpRzx3yQhPOz0cUWXASdJIHHmkEugVZNvEDACt9w4UX4Fw92StHySm1sml1fNON3wFXfhNKj6YQX
xAYo3QQNp4qm7RBYvSwLOznqQcZLJ0mc0Dkv64UenrzZkMjBYlUOcKsqUxix5wmOXwrUJAN6gz06
7yIedeyF2zlhJn7a/Hqy8aFeUf39/zfzSxHVvctExZg76JH/CHn9FtM50fCLi1YpbOUmfm1pdkfH
9D+ymrtmKzPkb7jYYStg1HxI+h1OdvWBAGs7LU1wgeawlzde5zuRfJqHdy4kXjSjrQ2KC/u9Vy7s
kHLVX5XqbthZMRsvo4aBbrIqEWWPWp4zSnTgVofNN540kUAvqp0WfASzalyE+Kxv9TbeSNdvUYLA
obhAQMCaQpcMpOvKcd1YO1/IZ2WvwG3KqEjsecytVd9bnmmxGMzqpoVFMEGj66QkNWllr+76cpjI
ukA3r3Fk3snzuclmXjPSeL3B73XiYoeusZl2DGdd9GmNq1jZNxaGyLvr5ryahFsT6831V8ZcCM6p
+GmsIJg48q7BLe6mS+7osEDzNyGoHfYBoB3g10XEt9o0L58PE6kuoD/j4K5BjdnB0Ees+fc983my
Gy/M5QtZBywi/Oz+cLP1NCXUhXSJAU3+xUAnXedCNgMGD4Qb3LNsYERn/6MRsNnRzyPJWW6zoMiH
gGHdeJiACC71EUAwpUa3LDF+yVMrIaH9v+EjliwIu3AgXQO60gbxakEMPQB7eipb9HRCwDJawr17
1pzGgUkHUnNdzbX/GXZzG4DUqG5GjYryhxHNhpOd1nlTAOAIE1A5kmeqqqHNT7FNoL2B7A2wcKwi
6HVbBQlkOyCotUpFy0KW+FBnZA7atRgjGeg97MPqy0E0mkvcwkh7mohbat1eT1U9jUZMpz2BFscF
AnobwmkWacECILG1AmdC4RhLZbas0Kh3WwRnDsEZaMGOetr+5Ga5uUt5izFRYpaZq/1qBc8LjKe6
ecsndcSU/AhY129TzMVGc6RMqzsmsdcWgbTXrA3QyMSuTt5xZKx4WhVdQ6og6JtOIAWjGAazfkEo
R84y72EKvn09cnugYWoUd6A1PJB8xcRFLS+Wa2pfYe9wwz20rXuxKSGslbztPJmGb6Rxp2P8hbpk
PfYpOgHQb6yq0aODkn9oPx78GvEobHl9o19nBPGhmWSEXRqmKhEzo3XnFsr/OGRqsnGKyfjO3Mr8
0ZcGHD2k22cuOKtE30I66ok9rMWTI/drGhxBwtRhkcD8bkd6m82/N7d/ZQ+9l4Zz8Dek074fbmhC
qA9g1x//MfDLa3Svv73jaADHZ6M1A2JmYVgq+0cmie3bqfaUbee8E6izSpnyvxSOpQGrToc7CvU/
+rKGw368yVM/pXDwTYKpAEAy8zHObyidQw3xatxY859puF6BabC3zqEzL8OI1viYjkGdoZUJ51EU
U2Lc/uT8VZTQxMnlY+k9Vs/kdwyOrKUGswDGNg9j6VybhnYGjQcIeI3M4lFurGNjajEbRoupLdXC
Z7gzs3Je0zdweMwBc0fOUG9SPiYFc4ECJ9S3tROTxiIV+w9VX7EO+l2NdYs9cYj+uFbOKsEpEQmm
+Um42nOusn/+QuwxCzfAjo064zkjkvsA8rnzJo+VwcOxelzxsAy59ecd6QAjVbO1ulpf/3ZdQQFw
3Buxf+8v5JYnsxSfZqNVTnza6JJvC/JVlSw9shjCJmW6hLisL6AvDg1kiNJZzQLKEUIElebJzJVJ
AS5kGXbgvCsf1j/KeMLvY0XEgW1/NfjkEsvFWK+UQEbuOXBxuQkOOOFLCGt9KQSMO/3kJgzRYgg5
jPvqmoEcXiYN+iiNMOfnrp9wUSwnJwd3p5V8QHWO/Ja26VwZa4/sM2ziMmCjIahclZULTzBUzhWo
qJ2tqPUQS3XPTVppst3ymupF5eY8KS3hrdJW0nl0YsocxA7jORulrXLH52D3N3GQR30H1iN3Lqv6
ZAAAfodYscYw6uaVCoHbmsCrVHXUESl7QL+E88NwGIlZ/9l5Fx8KzxP51kEjVtoN9GSC1yz0mzbF
Wal49ozxmFbBO5XtDoUFHA2pE6hHdE+j8887MEZ7ZHobF6eN0B6JUkSOP9Ai3fNfAEZ7J6DbJXuj
Nbdlyzr0RTGWILE/jyStrDvL3n8/P1NCiTRj1fmSuA5EwiIX2PrTkDl7tBEsixhjB4mZLeF/rtcU
LCIC35P0FsD2/d/26V76vW5Wj5KsAsNf0aw36v1W4stApViOnCvEGjDZA97pQ3wYQOdkivawygU1
meAJUy+MBuM+Tk+3FhkkUaD68g+2XMZRmJxEwSPYQDjYBLY9fWzRkZFYCzFsqofM7ok/Vab/37jW
Wh651JgxsMrYOw5a0LqDBHuhhAfSWX07Rw0moWrpw0C5dnhbl3mm5r4PzUvDIXJHy93lB8UNVEYQ
lCFFSx2PQUdJ+6gIzpdw3Jno9Tf2b5yzL/TuBRE1uCnHvoUddZcKIQZGjgV9zLWZMt1CxLIZ2tjG
/Qgzzi25SQ/tx+7OZWi1En3jGIpdSDXKtrkq5gubk2WXq0z+7BMYmTY4lRs9gR1ASDz5qTTR7Vyj
r15+3vrKEsGQXLpKegzXkbLBrdoFHNvqpSHUQThrKbhPEAXimtWf3hjnAZ6PyJdUmJw+ocrmvoGH
kKtzMJuELYIwnhDtTGtiAdoOjphVZils+cSAmhhLfhT8SBSbUGmknsQYQNOkC4nPccS7U+YwW968
j/zebeqU7E/pNaw4litydPD7DdIvutQXAxWLuLIYpBtDMksG5x1z4+ZPH0MY/eu66p7ZjxW6SN6w
5EowdDT6r1xIY/skMfmI54Gyy+qgoc9hRTIjE6CFnVQluUxwZCUGQWMLD6N9F/YfE0FGzMahhBaw
mNDTOfjyMz4m+mVX/jKN2Yh/wXEbZwgXGFmjLQPKrTeo5F65O9k+Mlrwp8sQBOl3DoV1zMB2mtRM
59xL8wrBOkDI1XWMBNRYpzbUnUD7s31j8/8G1ges/a390yQ2mkJl2C+2WIs/J6YYtyHgi5ET7HO9
luLHvB35Y7ETjdGdbLcif7Ez85+F97fvtpHma2yrsqt1N54iJowPKkmOnRxG9BQpOd52Hk8b4ZrV
bpVa5qgtxEqIyNPSm9cKNeah3cjif/pookctq9vtMqqMZI29wEiqzQwNNVGampNHeHNs6oXU0gIJ
V/Mp8hDQh53zAFRq2C7MdhI1Rn8urX1UE8LYzuYSb8GoZzcQdF8wGc1/0ddVREzMw3ibOfPQYThk
J7/3IZI9Oq8ExD0D6SQth8E4/zKaJGsMUtuonROKpaw4+DMjrKKRvuBJDYBbuB4IGcEc+Nj+LOGg
BLf0m+yQVC4gXVwqRI4yCqkf6a1JD9CPpLiUsMI3GcfZk4UjjUcuxLmAB3rhYn8CR6s3P8BeO22+
iEYzJ/XwXZKNcOD2u4TFL+oBbYXF30H917nDuKYF3PON7nKDIVfeVsfoyg4PDqhgeY+enWPi/yUZ
1Z8CuXtAY+4jWi8fhh9lYaEfk+lGG/1OnaQQlPr37nH8vVekrYTs0YIadQGy/LjiZlm6WpNPkhCp
ZsLJ4CaNuNlXuofGi6fk2PO7gKTJsQA8VoO/F0JB1iJOD5VNIIkCvEv5afBD0RzNiZ86fRsE/5UN
726EWwVM7re+t3moCS0vJ74fknUb6Cax1TWeG/BebxftO92fJGqBx5N3zgIhVYHrCS6qfAy5q7D0
8MNaNdnZX+vRbYTUGo9+wbbp+hhIKZGKwxQzLWE4e/dJfsc1Kyw7Dt/Kywp9nEhfJ9yj5vEu8MZM
zTZ5qun6vF1rxD4JXPEJwNTDBjt+CP31u6+61SM8PBakfVN+2FVgjhBzIfWwXoi+p9G6bFTfyz+a
/Snd8hs3Fa2QX9MApX8fyBjZgXoTtLU3H1LhAiJHU8Y7kFqZPLHy+W6zxAfLnmdl36sB/jXOE7lA
c4hgue1rUS+IhknYpIyXEWp5WLlJhJnfgrwmwcHLzKE9WkI4732Xi0h65svDZeo0OFKsi22dFT0B
5mfsDEfa1hUs/0D1z9e0R6KqjUaomPmc4PqTpxM5KXHMLgR99zTJlObBxsW0P5YRd6DP9N59Wk/i
XBp0+8hUx6SCONBT6ncZnW3/lHJQRQOymwVxJ5FQKvhW0/GcvhQZG/SRbvaM/14JRKsvAYrQnRGR
UJz6XR8b4dYYv6bFzyNz6DmeCvEs/oky4LpPKNzO2Od2QmI8MX7nF1UyWNcEM9OywSCG15Ngs6cR
qqFeTKKCN7nIdaJ0bqcHCaf7ET0/G65u+1cI3SNjd766uuyCS2JMO4S9JFG9sKGWSg6GxtJWW05Q
ZXa1ZVyg9hP+GhMOeOYRByTpOOy0v1Lx5kl/1tfHuXKY0OJfYNpJeonWJW4DPpxOievdXEYPpxgb
81sO9gjbRivQ5hzF4nREsasxzoABcLzUgodmm8ijFnCp9hPeANbighkld2XoFn0RlXHRxiXr06VC
8AgfE4FHHh3VtvjTZK3lxJisZW6BtXpjE3c/nA3Ki4EU7crHWvhTNnn6HX6aK5gEx6LcXlxaMGoy
vzB7XN99YO9Z4pD093Z53rlOfsUM7Fpk996RDZj9ptB55WXA9/6xqFyCvS1zmpi+ClzEndHDBHtV
GDqA/6BzY5BN+yPSuZiOuZjMPS7VoIs3obG2xAKtvocxT3CG+lmXbHBQJ9SbEy+qdhSMAs/GDVBn
U5Gsb53viBAjj7ZIf3gAvvqOQbR8HdKoCA1m1c/tm6R0+srEy4ReYGlN2kJCLSaUXwOm4gknUxcX
gZbPAYXY5ckob1G6LQcqw6oV1oXM6log26c7XDkbfro6tqxtR6D+8khDnnRPmt5B2A1lAc5ZyZKE
otAkCczUmAFpA4/vtcP8WeXzFcBWt2fx7dFOWqPomz0kc63RU10vJ1uHkXHEhuX9QcReUbO4scz0
uPmKDV8nJeFfAn78JfmBZ6YjY7Maurs4dRjU7Yt0k9D6ue9Mg29LvoJISMnTDFB5InrR9ef+n3k1
bwI5RNFWcF9ePSoTOll0SLNrVpycQev4vbPxs/l0AMpVB6xHoOIqJr1e7DBZFRM1/F4I64OWDJOs
1rrv7K+8e5bjZloavkF8EvkvrDOLJgoC+E0g4MXcUmhRTIx22qgcsDGhCo7t6vVSCYcaB3mEfiBb
mbQ8EiVnS799ZTzJEo0MykGXjB9UKtNjQxghZrlGzsTFrPWYBeol1/7BbyKcsWirHTPLjfHBJ5Kk
7+RmXud3pb4zx7Ww0Wsz0LIRDBSZx9/UbHde6XzCSFmUuLAVLD5ccf9N8P0yNd2Nc/8blC2GCCcX
aZumvbzaec5UkRA0GxZLJBkztVejH8qbRL6ilOzX9CGCZ0cxIm8NoW8HGeC2akB1J2jX9EGTNsVB
acGu1JxUWcQ05ORWCFFgxvjltshq3QnLOvHBo7qSG23ToJK2RvbgnzAr6eUodmEK9Ly0vHt+i96z
hBjhZVYZN/mOuiHdHCjejgwT9AtFVNpLhMg62gEyafiT4Re3p6JC9i4j4ixiD6qphgFJVMvKSFUC
0WepsIWythQrvcc/UxNdE9MqPxU29Jerubzv85yA0ZibaMNWNCLbxi/e+5WHxz3jC+CItZZaF7Mi
0/kYpd4PFz8pMQemxII9OnSA5bbaJ8eN9aH87OHV/S54CIfohZKHy+TPJXka+7fm4+mYAqA1ApfH
YkW4kIpzG6jABEGxw3N/oEdcCHbZhv1SyWW/SQGNyuSonIdtMYmPbxRkV2K1YPnOoRU1Rwh7sUry
lfyy79/M9/ljAo8wpHFkV4aEwDTnJ0y6TjQ3bBCADYPdRzdYup9BppzI9iwvRVgBFYX2Jmsd88eQ
YBsO6kXAAK355TOt1ZdVkRejqLvyc5jHoOBy1CAkMpW92XraZSq98uMO/X5pVI+FDEJ4Bw52HGZV
qsza1etaHR3lTM3t7oeDpCKeAiR+WFwtMGRK/HKvSgQ9qvep3KbgHP6St+WToBJ8XZ1cyXV8Lu14
ABSQNMLAjBrZfK8upKB85a/0Mb5W3SPXGpz/3NJVfsUtCGKXYzNmQiH42y7sBIPIRkk08RunOG71
Ru+95+D9RRPybNVeLwGUfvlf03sdv8IIIXatxQ6jsM13VnYJLOrXUUW94QYwi8k9K69eYe6Uokoe
0v23npdcnbJLSq1bUr3UJp1T/QgIu2nLGw8UGKzx5o7KJeAKZlK9WYguAP6sLLMy35txSKvw9wYX
wln+eeOPihGo7wADBm440ARdDgd1WMQxrmJEFOOqtX3DnDKa6lq5HFnxX3QM/kAYiiz6qi7grIN2
JTv93m+E9TFCnB2JpzJ/U7wSmNVEfy/dD6tg2BCp2J8Dv5D0bZJRzFKCBh2VDIYzErMrxuWz0mmW
h4vNQOG9XiO/w083bMLRd/xcyhQuXDwOlRK4fWoETVGgYil5mGydhMXGbs6vZI4muG/qr+Ad3Iv+
tOKK6mj3WSGoEy+JtzqfUqKkEKoJDqvox8ObovzNJy7MIaQ9utM9F2ygeWgaFBpYa0gS24KcepSO
ZYivq+W1m+2mqQN7dMxboCl1Fy8GwzFWoW6sk0xU7waYqoXEU+LbkZm1/HTiNM3PwymdVkArKUev
jAsFDJPB0fNLGZ0/NrIevDt4JpxOYrBBtTkeF+oeBYKg54bYXwIcP1muU0Qb03VA6sKHziTula2K
91+PNb4K6cnVPzEXApdLlQNTNkgUzRmrkVots/Q8ZVHY4i8sMRq9F4p9n+n81WQbFJlCkhxN+WLa
e2ThbeO2a65Ty+9O5fg0QLGdinpquV+Pb95Aui01E9T3EWJS03RRfhvLrbXiUxjnDb5U5H46VxKm
/OF8Y6gB4C9QTAwIwJTHSPb8+cA00viBzLf386tYkZScQbGwKtbXKg7tlPoRsPelpStUuxUcddQF
Z8bIsezKQoZrMTEl9HP1DCNJGFm2lJ3OiPTBf7ssPWP2ZXReiDDRjvzV10jBL3a+vYmfzExUVppZ
f78LP/cz88JrF8DdfQCIXHctImUqNRCVc/ErgmCxaRxMqpNhfIrhjXt4YGCHN4VfaPFE3PKBDpj6
n/fxmFB/Eq+2c+YQeosQDRM+MXEqwc1V0DWf2nMt5p+5kIcv08GNrkXswWziCXvk0yJECZzJm776
5c6lg+aplIFqBSXj8860T4RG21uN/tRKp8lsJTaVErpbX4nK9OC/wwMrz38gmaP7Xu/SNhQr6EqZ
h5Hwy/g5+A1MY4Lzzr7DSFZxUgzkFWfu4iZUoW5wwUvg5D9eobiknCfTsr6bvVwNmNTg8hZu1a28
Ct50QAFOCH1thH2a1pj2kZIQz3rp6Sga5julMNtS7sqs6howrEdv8t8W9cjEKtk7fV4G89C/JSWH
R8YX10YhVrFPqDFACgSEilVg2LT6hHFnaAVg92C3E/vlyszQa78v0x0WoLwWGwCnEz9LMqENVRQX
fCKZ97pIAZh+3L+1OwiysA49Xn5yi4dPrkqbRQq2vRpiJcobTBFxIkYaoLTF0YQHZFnNXrivEm09
hNht6/3FtkmFoz8V+SAzgdcIt/XAfWmqyebBbAqzWBqE0fxyFsmfR7E6BbJUQDc+XqREgpNIs2ti
Ipg8m9sbmxvsvJawQeDnsnxlv5doL26DrYda8JMDOGQsCKbrt/3/qH67m1FLs5Vw4hxzCL7ATsnc
c7C9mFHpSXOMaoPVYI8cEGD8o0D9DgGQJNxejz0a29V6H1gBBP2VHRtgRD60EfdNEKrmzw1AG7f4
VjPUqFWaDSBQs0V2YC2thEauke0zptAvjRT3OsjrJebWtBFMulN/Uaa5iQDQHol7Xu43tuTxKa+Z
Dd3OsNYFKMxQMbm+mWhTuIe0uI0jF6Zus6GX3D/aytsZxiY9Lj6w3MFwQgc/ZFrEBWiF7rQnaAIQ
6dSbpfCBN3b6FcYc5cRM23WvUuhB6SIvxV9zpGQtcMyBdicJ9PM4laO9d0P2yz8psXJsTU4+e6iq
FMrkz9Kq+58ucYPAtAJWEmkwGnVZOjSGR3ZZY/oI7RTuPRxSaT9BvQJ6aKHxkW+Trpjl1UmQ4c9s
uAhHZFD/ygIAqOf2wPsHB74KrWO9uatGFPZFfU/s8JceKBaq3Td0IOhbG438TjoH+x6tCRLmrFEw
ndwRouKAYYCnLpUAeSB+HG7XXNirtlnauYBNaAStOG1vDtsNgt3MgT9ueTeG08POVduFRp/DJnSM
kREf+swTHevUyCef7CV+kAafbpoV8CLczjrXSYYlWJUAsBp56I8DtYQUDQTrpKpMOjDiP6fk1aYI
mEQMLwkbQxoVTThDZpNBylOniBgu4XOT/RMtMjjjBsPiTGetTsr+SXs8P6ygdMB0lJY1bNtyEfF2
3m+gA4Bujjepvzn2SG9PNyXakrEudUj3hD3bKJhAzBI4gTBP/OAzCsZW4KS7Xci41z5/mAH8BO4D
4ThAZVow/kmJ+cYpqNpwxY66VirC0G5GDu5RG6GNZEguHrK7Pn4ctnRYxZItRiWyDRgQjTpbluNn
T5BBwsZQvD8HLhXiTQdWQFJ3XgM03tfxbDCGFm2LGTK6Tn/agHXRPgOQi8e6U+sC+r5vPnxx0Dq8
NvyLY9thoNv0dmG0P9Dk1cHZUliZS4ROaKgPwgodc4GfEbsPv57Il9p2y3DFgnfiEJPHBihweG2s
Zql/u81H6Hq0qU977OTnIDI6feRwH5wc8Q/ILrsEyBko/jy+HhKmiaDZTNv7sjpBLcz7nwwWnP/O
fpc56B6OCPEjNeBM/mhHa7Rz7L/F6FCK/UFVGGHW2UGggwYlq86Mni14R+Soyf+SPghxzLSCjbKw
nwhi9VbkInt+umjkSwj0S+wbrWAfrPqOZRq9pb7KqpRvBWD7Rxqvi0e9BhyoWnX/B75J+ZKtdn9g
tRp/iU45EZeVwIAwcTHsg8jVyp5NO3rsieLPjOoyLfuuOWzjANQS6CQdOGphaKuuQP9XGpFIQcsp
C66eYPYQIcG1hAOaL+Nz3NCEQUkwRun5zhdJiDXHCo8J8jyavTtJ5fkkeEF1iX7SrIFqZIQKffx1
TXMGOdU/I+8KBfxy/TiDSzK6mVnCckqFE49Jh8UWB3yHVmRaapLX109hfNFxVrkGFKrUVMONnjEe
rBZO8+T1Cdjv7/IV/sUO7LQY1yYKos7U/4ax+xBkXw2ATj2aiAMiTqseU17n0+RPDBL7Fj1+AERS
P8+ypDiQgn9jZ5ZfdQeRaVoM2PWl+QkkKnrYXcTCDEHChv+E7NFrx+J6Vs5pj9v16CwTsJdh5pp8
oFJ1GExye4iHXi9cUI3FLzQ4PBUNmviWw+bRcSQEThkw0u1fC6a3OWWddw/Z7U/rFFsJ3YloHGpo
L4fdSMp1VKkK6AUryoEM3Q7Lmmc80+OCDLPe+JPbubg8XZKxq8YKRExReK8+vvEUyfEdZeex12fo
sGjTh0vfb9jgPBFxYvFo2hqsN2GhcTqtattFb03B9PFQGHxoQGh1VQDqiEYhzBWHaKIrJyw7BWzS
2mKEtv1GdDMOlnOceaeNW2ItFLTHwaVgptNRI1Ne9msod3o115eDDHbS0Tvm6vi8SsYQH7x5n1T4
51QqHFH7DZrlNp37ANIIDXuTKAY7B4SfxiCAx7KlPBA6JLGThoyDbBzdHDr17gQ8JXPfgA/MJGMR
SnXm69dM2g0VA/kBGAsYOjPH6Au8cRuSfgDhLwVBt9RTlJpqKcHmUJfVtQFffKVAEd6Ln9eUBtAy
PGUkjvIpnDcyIF35PyxQv3s9G2E8nx/xSdNUeBw3HaJOgZlZ7R42416J4E0mzyPTcC4xdMZGRGyU
EnWGUsoeGmUyHsP/OrJYc1k5tSmi5EJYPh79af6dNlpB2/eD6c5NbaMA5j8pO/ZZ/F2GMRG2KNSW
8okKZFKYyBlzmN0uZ2JOWRffV+0vMTU1Bhrj0tNhWQiS7VEiMDd6qD4sx1VxplCgtde+wnswh5lM
wsQUsVYroZQcZLovl76gaKo18WkEIjIRAcIhGLI7XCfkw5imsGjLY3Du92efwdF0gleImD6gPP84
pybCZ7QPO4qEgY6geLYi9r8ayfuS2f00DVa5zw7cq9ZkE57S8brX2SwnXqnxl0KExMDFsLF9s6Yt
IcQ46Q/kAuXwZgXpXiPDc6O5nhkP/mwEGBxRbX1ggIao5bzfriidyVuUAr9TWSDY4aXwRwtAr5DG
vg7TxfvOePRBXmtb8ffpJbgwpREt1RiD7W8UZfuFVzeXrmK+1EMhwVyBdD6LDO1+LVGR8Imodko1
m8OsQ+TJ1Qhm2U0hTYS+QZjjDNHWiEXyRnFv6YOIe7QZSSq22/gtzCQZ7m6wD7f/mpaDjheqWm3q
whyfrB3Azs6SVPZSgVo/q3c8e3eJowHgndiaMW6b2rDpr09gK7voSNgSSpR26LqCh7KyvTeusyPf
bStkJBcAdDZF75OyBQpgq720cxTT31xRbXWPzzCsZtRFt3x3IflMW/dKx7JsaIpJOoI39DCgqqEd
uH6xe+uwS+pOX58FhS/DUHnacKxQKVgVmsBjLU3HU7XBR0VKFs9f+5ksmBSepxi+zznRvHOoNXrn
DqmEVSMmuymQy1A16stWD1cNR4oesukq3dVgBWmi5SQyMYu3fpHgElezNY4EZERv623oV1GrEj/M
tSMwqmUnSHKFILEYCTWwVt6o6ojVFGW+xJVDcUPmGxoQ21yDwu3dlk//s/ZFu2sVNWnU0FnNbuQb
S6XKoCvmWMgMYPsYhJcfpSD/xuE9VlJInnLsXgo8vdiQxAqdtrTqJp3q0SGLmwt1ZIH4NtGiOWvV
OeaPI1ZWyPokj89Kz+978ygJM2Bm/Tlk/Lt120rG5aXOYorMY7DESHXvQWlPHOg+5Kxs+Q12X2lI
/OjYc54IE6QeUQM7cAd9wmZERxm8RQiQxCjCz6nrvX0SECKbGVqYmaQW/5CwJG/kiBOQoJ4BJg7O
L1If5j7MxEtft/q0oWK9xLVz7gkv2oVHlSbs20b3CyATPQLUZZ62OmIsGWLVEvazLAawwHYUp9OH
p9nDQvnXw7XJ4GVjDqMkfcnndlrqXGAnWEpNcRzwe0qF2wD2ptCwIfZPzEkUPviX9GMSaMSe3n0G
l3snCUItFSyv1PVB851qTK8qNOfCNgUyDUOcyPtwl6j2O75Kl2StNbgkyY+ydbqGqUKvhwgrdZiZ
bV1BdvyoPe+j827XUORNrslHkhPnptwKjMy+34l5APpwyU86S2iIUUVqG/CdswUUAjmhxms6BSNK
vovULd/MsUmueUe1l0cLSFnwSk9e8VCPD0p7BygCyTrvtR9dh+I7Ef+B4opyiysqBMjb7Azu+gfG
VtXGbPgAsqtQUALK6MM5AhwURZRg7SFWy/yAkbpp+z5O1D9NFrolreH5bXwVM+uh3uO+jTg9u/Ut
w8drv5735LLjR4/RaUgVRGlqiSaimZSDtXJ6yp9ZYrmAyafPzUdI23QB0dOq9Y1UOz6zB2OMRBqh
/HSHsvstKkhrpQKb91tw8dk1uQfD/FpxvRR5ToWcEEIFcK6vbhRmzEnfyGRmG5WyFWIa0wtlQd3o
47SBS6xep4axXDvxwKz+rOSp6dPFQT6ayv91s7S6L2DZG8pKhF2YOoCczH2mwEOHCReCZI9UUY5y
RgYzydCxm6KE3+f7Jt17Dl6PS/0aQ2FWAj5Vy/jFcE4moLWWY2NrFCNSq7+TjwkvDTNuMdwLNElP
D72YvCE6ldZpVnnijG6zJVmP0uxAy24TnVN+L/6vQgHV51t1kF4i4csGjn1nLK0500dCXIwB381v
fveDnGl/Gqvy68e8Dls856QmdmHoWzfCd1tbfk4Cyc7f6Reexl4OYS7L5CTmQv3ueuo10WiSP6W+
oDDUYG6QFIS/7rMbrcJyAIiM10Bvjb33pGpvifK+erlIv29/fg5Rz3bo1deDBfmA0VCrYhX6ipjt
Vmxx2OwdXQfVXjP1i1rzeiDHDeThqqXxoLIdM+WMSsq8KkK4NFFYczaMdil+mFfI6K99sd8Nh1A0
3wX2Fqp+5iTKnWNaWjU1M8dhm5QVQJiZjNIMJqVbsKCZ1NfsLCsluJbBhVkqx3KGHh2kq1inNlgh
av122JOK6L+KPZxjUHroJiVPFfs61zqSR86dxZFmp/u+6B/quAQecCy1PFGiWtiyu5LEeYjUoIOP
BHD0nxAzL7AztR0xR3lz5cJnTXqgL+gv2Y4oov25IXdbCmHNnofextsRyqkcsqAIG7VpdW+pLo/0
ga7+dXgL6qCwNUyGiTZdZsuYcsY1t7KqgMsIGL6S1fPissAY9Sc3rGIJ0fJp+/a0xPYNoioD23gy
RrWXa1x7SnXoz4OATJb9VZkcrrFKLaDX/+RDORpJMXgQ+X+4CuwN13aX3gZRgQbR5XUtZ7r4ODAV
5Eopf+SOsYHiWOlfO+ks+GKlXMEkeW7z13nVlmSFwG2Mfp+2cYJTmHqwBSddlIhYQQgRmMeV6aZC
JL6DJhRzq/NgvPO8Zn/wbS/TwuY4p52dP8OQ7zAfL3KY0o+3adMPOhD7qPpDtzXUPm4kpKO2MLY6
dqiQ09MbE5B8G05b9ZDEPfl9qfxssNkBkK2xvquCnGNTqDmI1qtAZsZ/pb0PUJqgq9VVtPQye3n9
wj43IZC2o/HpwwgdP8DvgNeN1P77SxAv7dtoudKaZ6F659d3Gg5zwXucTi9wpD2pK0Sk7FFOCDwf
xzvv7YU7CQlp7XgLTKmzBVjLakdzeDONboM6XKLH6MrvvFhoV8m18BTTybrIYxU8e/8/0MtMrYpf
f11xNwmaVzCK/OO9q4Nyld0T3RsrXgi0sTWcBcEdxlFXrTkm5YfqFoz9jiYc2rHKsYB4cc1LLqgi
C6jSbU9SgEpQk5vdcN4zIJlbNNzlgFvmxODsCNFCuyvQwwWsWyReTgDk33kMMsZY9d4Eo1SgEjxx
U+mI25R4isWnMCItqrx/ritrG9oW9GzkllCfefcGGo8H9Bn6Ac6UAEkiaExoxO1Uf3bxvl9Q5RU2
9Dr4MzxybJQ2GDkJF2+eh1qLEJE5oINOIbo/LNoW4FzTdSXJAcUE3gwDloTT2AolFevilJxyU3R6
os4/fLhfiaCmt8B2K1mFzfpN2gvVci+z1OVKxTXPBJWl3lMDjtRAEmi95zfeDBKXv4P9fmlIKCIf
YJNfNlLktGahL2Ifx4FMLBV0wyA10JzvGGP+JFbJh3vhNgVAtIn7J5QFwCv8uxWrh/PaTU1p59Zh
pk3odnz5pxIZTOkUx++nQ8lD32AFpMFnaqXCw0F05AUQbcNu8Kf7lz34X3HqL5yw+TPuaz0XNJCm
4/BXLHe70FH5a1difI4kvgzO4a4vZ43iyZvHMDks5BLHQPLkyQz0kMPQHd8a/Bi2XCOCBHVbRbVs
alHSBaIScP3nhw19MJjngg0WxLuEzorNdm39PWVb1Idz82sHezr71Ucoyly/AJQboKvutowaw5Vp
x8LdA9yRS/x0LSSueXK9GuIVnMpDLE+xwDKngUcSHeI+bWRXULsWO0WA60ud8xiKCJZcpvIvZtKB
SE7tTCojJh7vTtfKGWAsKv5TZz00Bq8R9iEay0amkuQw6EvUMhdTp69cVWlsrh6zRY2JHAhf4GcK
h/ad+uJH3u2ouY7rurwI6R+aiSV1TQJiSoAhklIIyBzfv4hUDAFBqF6UR2dY3qnbwJEvijRiz0Hb
zWFVKaKDf+KWHjIV/frRi6nPOQZPlmxa0v8ne8PWcXQHfnz9v2RQDJuGilRUe/+1qkJexSBsuqLL
mGd2W1lfJ7+/DjFbi0LkwBGHJFczpaqEmQAPG1tGg7tXoF1+Z5hN1tSaNuyat6yBCSQC153+9knZ
EqzS1JKIln8/PpIya/q8oQy548e32vy0irR+tp/SK6vGtTjNf0sWnPPPNvmrtfDqhnj8hOm9abY9
5Bdgz0hkR2Fn7Wq/P/uuJ85gK2DmajZd3uITM0gkH/u/pZIHIoJCo/x/xbDWyyXUR9lCAoZsIOhQ
HgWGIM3zCsY4PzV4v4nvcrpQlfsfPlIWF2rkUW4ry+HC/fVIYiTYXLI9HAvJHJ+NQzKNxTaK6YyQ
iGvnip9S5RB46pGb9O1dRb0+1+YqPsdM+DDKXvvyk+X2ETbr4mSygqorXa0Z4zxcWwuPJ6phNT7l
sJbNp2k4wXD7LtpOwFtbXZseX251euC1YSY9o2G/SZZlUShVNMcCO7A+fZVTLFs/WMQ2TWveQAxD
psl6SKqqF0el9RR8soQuQj4TwCQ34j86jyMFOMpAFi/g1Z73Xbsxeu49icLkU4SPVp0yOccMSh5n
4k0XuJrL6ZueXMC4zMfjqBao91MI//PHoxjbeWg3rILDslQrY4VXgiA7GjS/MkkO/ChoMghXLf2N
5SX+q9RU3mtu6JfPV4NYumDUzeVMHjnFUugm1IfEUSwDr9Tuo7Ug4sq+PK/dDuUDCdbu61biHZSF
Rpe0Ppd0387y//Wb9qMHadaL30UQzSvxsP78W8NXl9I/XSSO8jpg4reNH6arJ+WrngviqUUXtAOg
Jk9PnZPFTs+wDdvU3UJeoqgMnj3/NEheld4VCRqRXzSBX69be/6/mu3XOO+Z46USyTVmaJmE55tD
floylL19sXrQ8syFETG4CDatuIQyUVF3aSwf+SkkMBS3PjakgPZDB4uqn+2n1Q/oJZ4Jhcenzbno
7e1VWY43u4czXyAoPuDLSxC5LeZVls1wpM4ki2WkHm6xsE3XcdgL9ZxmCjuuV7nwpRVkun1/mF13
rN3KAsMYkLIduQ5qPnpm//ntf/8lCW8lB4ZOv8XpC5gAVx/AvpNUhmxdR7Xbgw7M+e2y4QZC2nOR
eoZfNZvpo6R1tPINZ7vFarBGBxgRLsC2dfREVzU66z5No1J3ly1j/UFX223fYQF1hIWLPKkNWzzQ
l0voJ4j1S0dS90/Jujet1YOBFCS8QRK1ZlU9V1BBKDttrlmZf+H3Q6491W2jmMRZHaKrDiiBFxwM
C0uuipSHUXAIHLFwzxfOoAVO024Vm/sy3nR23lWbsl/s/V7VDg6SL+6QEQas3di70B76K07dGw+h
OpUGCocQ/3BG/78sYKf6z4tWbLZrw517Qk0T99LwPUhNPXDOAVSr+LkVqU0bKMAyMTQRjf9iuuHu
MxirTnUMbbxPkxDVHcBuMwEYQSLpNb35gRFL6f5YKyyG10Xu0W1wyqFaUyb6KUtJMGXLr+gCkwZF
xol9wj+ayPOIhFAYy4RWNkq1fqYYZp+fXrZmpbuQOKbm8OiN23mvHuq+x0POxedSS4QCkDBSM/Xz
V9JINROKdqXo3Er+2K9kyNaPvmkWxlKqvkmTwwrDGJZGMm24YO6aZXa5LytszexkfO00jMbRF/N5
RmmIHiSQtyx6+8c3ejDhgWjkBtCNBsIM6KUsSGvw26d7DFGXlyet2EGn9dJry+g4Tu7QDTHrpDof
YHkaiufYFj3AlsV4wo5sI9DXc1dVWHeYAo9TgRur00GfwGGZQ0nDRV+kVO72aDN5zq7cKedGMVQx
u9lGFfMxnLC7uHsTXH4S8MTHjr76UBVxn3YwWKSBkca180z3F2jZq8/oySc+TTRHudbcQAJm+1SA
ifycUHqGOEcJhX8JREfph8QW+jeqlK5uy2tWEsVky1TiVCOx9Lkw44BOo642ky6W8g64cnhMTK3K
03I9nGTYjOhMZf0j841m4OjOEK8QAwJWO65ZMLMCgh5lH6HMKY011Oi0LMztTdAVFtEZkO8UfFxb
kH4J6SX+h4qtNQs3aCwA84npM44a/Dz1lefRbDK91A2q6NCOMMfuItdtXnYF0xZN6VPZLLU1Tsdv
JvDAS+6wVYYleQPMmlg/15gBrE++UHEnSY7V09h9Ojb7Sj5Qh/lhaADADVYfMTjaSTeLbRZdTuF3
9G8XHiCEmlCJ4t6ztUCZ26eyziWz2QsmEuZRNUJ+tgQCJg/oZyhO4hwbHU1Qa1zWY2b2P5TLYAgj
lgOnc1nb+ePanB7yaDt6ILxVtyjR+qAwTPXnhDx1NJvW6vVTQ/Mvrs06SjSrxvrGOrxiLcFYlW9w
jhD9/xBNXfwqXzFY3tCs7WWMqkw44pKu1k4wzEmixaw5mTuMZPRSBMHMwpaOY38RqrrT/dmdCySy
t1tcQg6EdWvFHY5R/U9o8N7TFNS/SoQAxaYy13TEghRx3tJft8nIf1Gq1rTEBcsQFUIMgA69mT8U
CLVTDIEQIWtqWWMsB8J7sRjrESnWEcY/ZfJCqe6DfQMqSgZjy7OO8HOlQt0N6qu1zrgBJkn/Z/zm
BR6kkaUbkVB9IrLf8Gefoik4I/siXXZDzoT+sasWSmV22QS6ytHy2YGCAJvB9xh6MXDFCLkBGAzb
rk346SLtzgsVHGlZ6wI9f/IBN04HTdtun5BR3CKxL+eRCeuWUbOJOh8dJ999wTVLClzCGgTnnDrs
xGLRN9jyM2HmRCTyXBM1b/czJvM/OJc2+QMvlwfsSOJbmDAvUkFDXAimXNIIeQ6G+vNzKsq0twkC
LWciVeu4dIOCEw48NTTnnnW2mVb+fGAJuedDD+mS1UhtzccT5m9DkhXZC7X+MRlMfjW12Gn93awL
ETlzdwgqapbyZ/Bb6YH43ogg8uoci48jvqtoLB7Qv+PGzRrRNLZqOPS2k/bsNN+2EoT4p+4yxBdE
pZz6OrHL0zuv3thK7DwJXQ4OIOpDPHP89vh0dZh2eotVdRQt3xDl0ZyMl219VuS1Y3L9BaxzO8oP
plyKX86qI01C+pDnljdWsJnPWd5EIo7qRX05kKCI1avmSH7mla8pA7CnSlNrTvpZ8800CTsMf2Xf
D2PbX22tz4FNEnlI9YbVL5Ce44E0PMQClqyArEOmXRD3HHGXs1orzoCYpBEnZAxw+x8/FI3VlOuA
AWz9UhSaWk/UFQ6PMp2Fc28qf0GYtT61rqcSvlxEImX2XYcqBOZH8VmbldHYPVFZ0FAU1z1E5KKO
J0asgDvDDNrHxPMcskEWO5Z+ElHaxDJlwJ/Yjghq5Ts3CiEeHlXwfrq8zVyituKpBO2bCiFYMuyR
PcxWzH3ChuikXg7wwjM7coybS+ebXgIGubK5imUAa7BRazmFGFR7UACXCrTLO88bO/Qs+6gkVe6O
sLTIqyK59AnL55TmucGb0R/evpu+lv8yHv6CruZcx0o0IlTNfH0uPl5taNg5ymbD752XtdH15+09
bESNdXDLciy1+QQGbtA2I5Ar7FeU7M1bEqFWq35H1Pxdi7NyUibQcvpXKz4TL1mxF1zjAxy+ug33
+/4H9NFPCfvR7+ohLfZqbcBghTCEeS1bPR5J7FbU1QIA7E20vgkfpVeasHToI+5dIXxR8TtAmh+q
9d7CCIZyMGXSs8RK4Zesl32plIfndktLI39o6aBTH3rhHz4h/BLRMMib29Tj+SLygGPVwBHRrjE8
yMKC1cnHAVgUzS0exqGXc1pk+DmVE5O4kHRLcvmEdAPIRMA50i/iT+rnbIARHTrVkziYzIFN8uWE
YGeIT5kf1QQ/P37C+nxH5jV1w03FFStr4T3uNDFyyizFXWZZJZJ/hLXlR69k/RcbKgZ4tbcr9+0r
s6e2SaoxO/f2KB4zs7QNOL0xQOz9dXQQrLZTgead35us2k6ZpcyqfCUvQy+o+v5UnYqaQedTs3Nv
HfZTTed1+AxBkuXblcS3OlFotxQT27OSUCd3+yEGClITLMuKjUSJWujIi4ARy6JwuVwoZqlBZ1uR
CBP0t5ApTm8h4mywkd6cpfc8e+K1JgvgD5AsVOxT46ww7FCq1EkKkJYDHGNNzVAP/1mLT39bZEL3
JwaaEAFMNR1TnE9vkmERfbQar+Xj5698X+Xx/krK3/drFRAjnCyZWCC+1Q1J/v68AngAnia/KUGY
isdEemngvawM6l1OaiE3zLdrtmlAj/r5RRHeonv+MqfvPrwycG2fJXEvmpL2X7NV+HEayNl0+ZrX
3B21XX4ZU7z3uSrkOkVGj5YVwIxzJgg1/4jg06JActMHNEX86aaGwLY/CEOxOx5w3SGqsxPe/Rl2
h5c6brNPptqUt6oWMDv4AMpZbqgGVpvLt9Sw0QwwSgg07tKBMMA8Ax5LzK56YKjAdZyUhfrEZR/3
IWNz+2Y/3bQLXT3QXMg4Du9Xh91p51+1IZPNrZTU26ylp42lu2XHaaxIaeuodL/2AxEz+UsZ7F5G
zirAqyp4xGTWzKGCyKsYxWCpAA2esf2U4osLpiKaCntngjeujprH6dqQ3kwTSirr1ztWRyNEH7rN
dU/Xeh5tG499L+xxHFvIYoIQ5IE7lr6uHyCHwTA3zX3HQ5AfB2L/FrKuXnNf4jLVg994sUOYdeIN
5GOykenKHdgHLvkK4o2Hi1DOM2HjRB1aLsiffMGeEqu6dvW1zTJnAB5YxpCTPnEzN4xn11ZIwHAT
wteevS2QWr5tk7P+oJrRamu+qyfj+EGM8b9gu4MQulupmHUDaOZEoPcUhMLnW+mdjjRvrhNN6hOU
b+xWOFIaDEiqPVk3i+R1Z8cS1tsmjc0gfRRxDthBm+cIoqpxyl7qQfHvxnu5yfsrIvYwoQt+Ce6Z
FURgkDuf09be49fHhLpaXSpy4v0Qs/PUaODa67Fhf4KxAeHC06eYa+A9m9X1bKHM5RoPBPBryujn
GV3+2NW7SjZbNt4x8M0PZMUbbSYJbgLn7ES/yt4VggSEyTTRqlpDT7KjDBYD12BeLARFofehluD8
WEKaFMy5EiAmol0gEM+hMH0dGhVozMqVSnyijYY7gZvazqfUekSGZmGtGxFjWEijnH4hPgqdMizz
FpglRLUZEQwvPDTxOgE+fKX9MGx+GRyPyLbf+5WWLXnTFXTFkc1oJfbdEqP+2oKz0N9I725rSTBn
rh+6QW+1pki6miTlb6uFyX+Ao8e2FyRV+Gt0YR1p8BYfspbzqkZK6RJqCHR71XJIsqqpZ8ZMHdyU
LZElfs8FYjwecb1nWJ01Afzpt1BwCitl+T7nK4lYz7xDaclOUwUgnpO5YS7yE+SsewwIuLCwyNOa
TlDvBXnHslwZxmHgDtotnhD3T1A2teBqPKllHlK55oYw9POio25EjznEs7LHGnA229yxeq3qr55f
tZb/1mT62o2ge5hRi9fSYMsClPCjh/OngYoEUQxqBO1/b4KMdtkgRU/+EgEGcsVbblFUv2L6UHbB
G33AOeGd4/Vo9owixfVqnGo8wXBmY+IQnNoeefdYnY/xXSTzG1k8E9y2VScKEdW3VujYCKcOU9rc
GzsJcRXYtU6IpuGat0P4aMjhPhlfl44OeMwDYGeKTC2eOHVkPbpnJGh3jBaQ10TEJbC3M4w5zY1F
DpX9Zo2qpUA+TvHd1GPAHzL5I66SxmgltEJxYBAVdp16UcGFgUKFdOx580OeMZrQBOrteNs92Uga
VjNvPpZbZDtTxyOHcukH3x42TdrUf92BNZJbHBgYC/d7513wIolqZN780dbgndIswGb1rbvywLIZ
aBAoGXkIEXs3Uefq2Hzg0rKz9mBmxYk2yEB/k8IKYKp/eEFOCUwUUoNpph+MC6zSnWuRrVOtVfat
P1J7kBjVLfJQeTPPWfBglSXNXfwjQp9hhHsC19QgOWmhlPuqwIJcAn5rqajkbbMqH2xDlUjKFr9S
ZT4B40u8ZH7k3XZyRfuKDsC3RC7zVoT9vFcOmfyelGeZxVh491D7+mY6rJHqEM/q/Q2f5wgoqRHK
5bkhjyU6cqZNP/wdlTm/mW+Z+YpWqRr+NG4EaU50meZNcjzQqvaG/wTVEle+19Nfss18+LxWvJ41
Px39mIDcNIe8HZFtYndrdy3kuvbjbkSG+rSNPEGb2H0G9TnvmWQPnj+vzw+YWvtoGPwB+E8+XBRr
1vnrcL6ro7/lKXUd1YPRTyTmQ+gX00PEWPTZRNCnoo58xeSoZm9K9Q8IJM6xC1y1t50p+9S9O9ti
0AgEzLZ09iismwcdXJvZ05EBWtIhs5yMy6yfLPzQuYUoTv57FIe7BxqvkWGn5HHEzU5yuEvc7kVE
wUjJTh9rhV4cMADJ/CteCP+fA5fSc+VUdNqLB7sPMZu/o15pF86XnJQoatBI99MRUUhxwZtfPjOZ
zUCA33d5y7O2lw45x6piIuSEs6FmsrBpsnwBJ0xLrn9eGP4W9QFcTWd7SmQpyRdF5Quo/RLdbFxC
1ECT3fMRCZ6bqWQKfXIfwf7nqwJevF6//aFXtj1rkDagJVfl8wLV+BKjPibTm7Eg0ywCG6FaPUO+
CyrJXITJh+jxVyYsXiFgmxmwaw97KFHbJuinXK3UGBw2mqUrxX24vWJT/l4mjEeP+zi8tv03RVWa
FtiYyjgXHxxP8m+i13FThDDxuCAd9sHyFSia4N1dOFPrGD5MSlg1iwfx7PKcwWyUYEqnrROkAJTS
j9gchBQ8Zmuw4flpuVn+GW1s0K20ASRvqeTORne5g71flmHSNhVLSwwUJc6bokj652xsbR/zvevS
LFueKc5ApMJwlx5qVeIVLJOb0ZRz+mDeT4QiH8rNOjiSiiaq6hE40axRKy8sz/+Hx9o+S+N8Vz8M
TME0meXeh0/xGAnNz4DhOeHWWMLSgbjyOY6g7AuxUe1Dzf48AHmlVmJBkC8Pdl6xtIbMfezBEwBO
9ruvcscoPZMBodD1LRCm2Wkcahuer3p06rr15kKPcG6DOkbP+fiViljLarpji8q/NlEhoElA44pB
XgubHcYGXdsZh+WrWYIMLVr9AXVtP1U3PwbP1aKRWyIE1bUEiRA8dGIIXIvWc4WYozOYbbJsNeNq
Npn7yTx/R5RncD31RM2Ce8tU+ZaC5tmRsskXSq26apxA0/C6wmk3gTYgWMXP3+a1iBAV2eYXQPaS
XBbjI4V+HTixrDIam7UqYzWDjMNSQ1KKi9KWtSNO6MKNY5U+nXxyUo2lYCUTAz20kYOuwviHtuvd
bLBMySpfWIYcSbZTWsnoVcBXgHWFOSC9XpnLHLzURqbrjLkvpcH+VAQW7dhgC47SNd9cTQvOXZ5l
rKvSEv57Y1SpRPTCEHBdYv55l8BED/SZoPBzFGCLOYOvl+KXGJ2LEOuvdB+olllPIIgWLGvY2KOC
BNLdZZxUKCQZjzHtoh0oFhKlDG/1EQQ7ZW263Xs42tBkYGz83kmzXtNlN1vc0yk7GTitGPm2QFEO
C0GpHwVYkxyqS9LFqR5/Py2vr91Iu6jallB2qob5dUjxQBDsmNfSoxmNSP/+c+bmyqe/dm1kn+pc
pCYwDLenwpahomI8IVhOQ8Ef8MIl1PHphnw+RfUVFe2dng80t+DVgDeWb2h3EfI8Q9f8Hs5WnUHK
4Kz26uP+lg/vxEbULaLTZ41EdXZfMqwqP8Dt3OKdmRId4hfaGe+kwsINk33Od3SB0N+jucP/C72c
k6G+MpY1IsHVtKi7Hr7LWx92/pqIzfyB/qEeCF7s2/HHbnx9ly5ZCjzuJyeMiGmooG9XJA8n8e+d
JmZvepxGmz4Tj3ZRjyBe/DsS0ibAqVhf07c0yAcdeOT+gRj/4xr6Py93ltykGHisYhHC6NC/4Hf1
YvOfrlTj07cg1ILXh0t4L2TWYoM2N1cRw0HUSz/TT1o+Od9livvfFcSEYDD9gHMcrhVJ5eisZWXy
sEcayXjO/QC3Why2A1lFvvM5QmC3zwrf/KNUKSOBIQr3R9tZjoRdK7TCSXO8m8uNBTa+Qpj5LgIw
YIRxvluEL9wyB1VHSkmFFJOQE+ox7nvMTOGuxkg9fkHMknTBCP2iTjDsXmZ7htXOcUC5UMEbPWFE
gCOIlHiqughlsoWJ5VBZy298KPeKgC/nXz7Dmi1lW4WbbnzP4kgDaseBZ6fYPqno/oaL/hJZQ1+0
yUhgSVo8mCS1HFRDUwgappNYquCw+L6TM6nt2Ijp3UTKalrYQsAVA5mstxd+mQp665GfOo11OugP
/7bgK8kh+s3U1/nr2GCKNVN1gIB/6NB3hVw7s3wytDrukl5KfgsVv21wer3Ra/95FLdF5dyk4bQd
asO8prJv8WmQpTDjTnmlXYOMc/5OjNChKa9BlWMhGGvNN5VSf+n3o9HeSGcJ5T7CeQGd0itsStGB
NjcKfWNoBrDRwLGtarTe7FVojca/Kf8rEGsXBySt6Qt7C11vQjvftlp9T77VEMdOY6GblDKWbjGP
NMW9xtmBaDVJNCJZruF7/j3CmWZIAXR/KJtN+TDW2BNctcAoohFh9aY/Wfmfyx2kT02g+k2XtR5Y
ufNioM5IdJnTb41LckRLGryZGy7ImmMEbB3AZhFeAG9e5D7fecK71vNhPc00GslUtsi1qqCwSf06
7DwOsNBNe5HeNdTXEXlh0B3bRBm9ZJfAFYGf3D67on05yzOlLu5Gth1FPEu14bE86WX7nNvkDkFC
7LOa5J9iKzsZS7Sw/LzXwIPuR0YQQ6DFhJQgDe+S+98INRB5UaU6Cf8qNosvG9BCLXL+1GIzmUAO
klJ2CrF4suCIHmISIt9q2ngd9hwYczu+sYvl0/M3kq9i9FulUs6U3AymmalheiY1OxXnqTaPHKml
AINgoUHHSQ7O6oHnP1HR1ZLjH6DBnVz6exNI2HmXI632PWBJD7w0Xm8Guq9aZdBCyUU+vL3R2LmN
YgFF3m+F1MqeUsFAzHrEOYENH31GUMvXPRa68VQWBFoDmQMfQwS2rx+VrPv8Lyv3B2rFOK6dxqjy
2GplAt/d3+Od0Q/yWpIbrhdmSZQMWeV293tOk5TV04wTpZ6OM3AyR0IZlheWPYavNsaDYIZxoKGq
v/Q7qtXlFQNT2wRmd5ZH7yL28HHJJM7z8qMt3X6N8OUyeaev8sA2gP5prGWGLZ6MB1m7JTm5IhGI
aoCwpRAWbYuOn+wMY5eKLSAOAsFpECkKV4J0RXIcfIkEFOqKhrJ4tyaOREONTml1JeaZKK81s2R+
L6tWXLkNM1ECwglkzb5NPdtvD4uwAU3BrXLIMvw3aUbGYMJ4+THR6Dw5tCYPgGBrZHMq50zHwmoN
XzwtyZbXSeWx9zeWG6Gs7LIUwTtODgt9OZznTsfPoySXrf8xDpsQYKJxuXeuWUFY1n4POqaiD0DP
S1KnlSatyFnGy6jUuv0xY8Z1m6EN4ypW+S5c4XWM5kyNvIBF/3dyqzZU8+lcOxsSMe0oOzFnikUC
Awq67fsem0c8pZkqBjQVg4PCCi0RANBVkpRqgqpGkR97M0Acez0GkZc1rIa98W90qPuR4YQ4FgVE
f41tO9XWuZLYAtMm9JwWg72No+NiIB1INUiZkIdW8b+U65S8EdFVQ+mXf/rkISF7G/5Ee06il0dO
+GFWZKVQVUkervpMpkYbcggxs5iqtdQcrlhFQSWNTAuuMZd0Py+QzWCZu5aVp6pPZIv/lu/rEIyt
5M3pYra2OHbRg32WhhXuqChn0/5FaUGbQpFE3a70MrbOi4Hk7pmVcroWR6SfVf6bX/LMmXlvXVhG
88EQdxdUqOT5eqT+AoRhbIqO64QZC0xXHI/wBAVb4CJ3dnL1iFTtXaTbwCjUzsXikPhmISmut22u
BMeVK9jCaMYhyo61hPmkdh8Lz7SSK+/16hjvya50c1p9KP9bIqQE+vDebpoaV9psmFRVfrqJMjos
rSgnkuAF1Av5D0j/rHkCFushM7jBWknxr+gLZ4F+iQ/glFop76qDRPT/TRuIpiEkUcsz0doTwzjA
8hKN5qTA/Dm2yEDAjceOt9aHseIPpsLt04byWQvYfRukVIjUM1bXzOpd9SVzYxnlPn7XR+1cOCRi
1Lz28s/6pIKpKOHw51wi8rfxNOgh0Uu5lwghe4UqAhh+Ja0tEd56pqWN5juJZnpFcrYw1OKtq+2J
ENnNpP76114jyizS5tuEtHSDKEqbfIR4MZs5wLuLfwspy0nnb7uO97QLM1qN8KVYsRmN1zvYZiSH
6fZX/UM5ZFrIPRe7XeOXpbMh0Jh/f7cjwVXQHvW4dvlBwQ02m1L924DODF6TPRcvNp29dqHkig2F
YAa4IyWwhAV8/oJERBpZV0nalvc9ETbcvzO64Jy4QGRh+SGGesDQrvea5JvQSvmDFV6Tv1QEHADA
cHcmi8QicGYxBxJjbQayeRNiALuldHoHEqDG9REJiJHakE/9mNpVV0QKEqZZqqOs07T8pTWE3VbE
m+hTIsDlGdgwEnzVgR6kSM8nw84Z/HMsFK6fDgx56aejvqyTopQbk1w5puCLeuui8kDwa7n5rMyq
6/oS24hSUfGYVhWXsTOEiFq4TBgAGMOdk4gAc0Nvv/Q8AczInVARsz6Hd3f/V+xXSPaoQmPABT8w
kkThvBQJQdGHpE9szsrtmOGZkswAGZkdTc6AeszCiMbGw40X+mp9FQw+dW4U5x4aMDmcMjJy2ON9
S5M0HJjLnSDSN3lU6Gta0oxJ97kLuq8nUVTZ6ONc5X/lJe+0wTg5nldTFmZqBgnghvJpUyR14uay
aeiDSe+xay9gI79NwVRjGuy9qj8fJ2PqlxzfN4O65CwCdhyuIetSpvNZlWrPKt7yNkNromJd6gGl
9vDtflO4lK54r5hkZyM/a3ll1Q6tJ2Q1KQo4YI4DK7UwsY8lQDhuZgg9Q2s1P2u2EEkgHwUCUKdm
ASwRdWj5cez4VQlchCJKaMTlFYmSLM3g8Okk5mOe/Iva6Ht2vflkyAjbU52x5rdNrM1UxgnrU719
787mpDUxhL1R4bjMWahBynqJu1AM9ndtfBgG78Jr6zvGRNpH/xUk2gV4BkMwZiMCYn4lp+8sEXiU
fIr4De398t2vmw7CNEzGjoeZ3nBYA/8BFbUlSqBbPi7ynlq3Rsx+6IRRYcDCtlC94N4JdQDCRq6x
X+2ZoXjiFy1KnIh+Vg0ffAiDHXQDGXijPgopBA7vxjV2Tm2sDkzIxim6isYuA71xemhphOYiKr9R
SUzJZ5Gn9jtFDjx9KAsNX5YH4u5hHuOaYFC3WEefpifO9oon9atcrZYllN2EFUMf1Pyo0R8qXKm9
ZwR5AMSrtc2civ9XDs/t550G+xghbFNZsqlmWDN/M8NoFl+dQ4oQ0EuscGzsnWKiBAkP/iRIyC8T
cQRKy5M5EaP63ngwt6IkGL/0asL3XAttdYvUDf3kTH7/TxYukBxW9/zs10Ocvr9nym9GpAl9VoOZ
/SWJ2S+9aGUgGxlyeY/DEaZ4X3yzREU4eTT/godefakRjvgYcnCd1Pp9AeK0ArJ0NQBmjIKER+DO
GPN9EGkndjJfMlBrZdizwH1E0feKTMM7hQPrD3hvMafCvx0ZDks9Hl2qMEanJX262pVv1SVLng2T
8HM4Kmwm3H09RKHBmpTkc2A6x1fCVRd/fxvz7CN5KFJxYfQdTkKwZi6hQ/tkopOTM50/WLGC+t55
PhFsyBRm/KD9nfu7FezIjPglGy8PXeJ78CkhGiRq8dnLstAWrmJDUx2HIjgwk0XRAWWHL+aAU+3M
2+AoVTFyxn2KKufy9H20Wf/Dwd2fnpXNZN6OpjRObY/RYnztBs3O80q1O3Cm4rs66ZWA8uEZS/Ns
Swgam1b5CZ3K2b3KUeeWrofiA6uuhAqNJ+PAqC+ZHzGhi1c+uCyh79vPSGoge8nL4UMbMqH6F580
KNbCigtsxW+5yhSfXzDms2Zgp3wYWu3lMzN666755z9MeXQlb1WdCDL1XRkYSmHqEv2bzYZCOFUx
iosbKiCmRXbXIsagIyMsJAAq7b4WCBhZ0CScniBW0lfgh+mrKefcrb0ESMkmYLC9xpfA2qJvGzVF
vCz/M6+KdXIjaWP9euY2zyUQckn4ciK2fXJTMktOBjTwBb2E1eUIg+r2sI04p6G3BcPsRO37PH12
/l7ir9UNodD73b4dKcnR+zYLlbpbGmeN0XCKmSl9ZCPEDAccfTiQPUWREfUXBvWK+pYgxO7i5xmL
rlnzzGTse/wlVLNLkbXgdd4nAgYc3/EtLC8e3DH3uzGjFWVjfWkKl2EeGSRf0Mqj8jvceXOiS7tC
pUoNdmTsz/gUfCF0csrlN3MuK5TfpCSGf1oVaneF3Z5+4JwwRWyJvqXr0KbYVGr+BgRRILXN4q1p
rGrZA18cxKwzMphqoQhxpcC+dgcxEOVIOH703anQ9MrtPfaX/P/WrYJYFELjXb0GP43a9CqKMvo1
Q0q/gFHyn34ltJnosTPiPIMZXhPr3EzWiNWXPEXuiIiu791lbxpccrSU4/imz+O511vpNXvrnwQT
UdnOt7KZoIMT8DRYz7LZMFteAYPQ+VWd+ieppPaWQk3exsaUD/j1/Zo29ReKL5+BdetFafq5EVD+
MiILLogEKkz72xACsRfEAWQbfCjnDMQMuFbvtv1xhO65BOIg1Dqeo37coDhH+l8h+AqeeOwcI13q
RBdAq80edsLc+C+uv2PIvOU5mXhyUzoIq6LDHT19EtU//5JzwY5tojj4SsjjlSVDK4UY3TwQj3de
GOKDoPbLbqPjZZFZBC5CA5vZXSMW9qNpWKlYskOUlzlW+SKyVSSBo7zzgsgU67vLM3o4Ge4n3p3X
XsGTm7mC+s0mtioaRd99KXf/6KqHGRJn3MYAfeu1N1QDT3yrtHqqwknwIWJ02cmPT8EBN0dWLjbn
YVsF8SBEN/mfTfgix5y2KaAr/iNLuy+1//ol8JESDKp7jmapJWlqfNQ9jQjVgm7W3uDptEquRkKA
WBGxlIfYjeO/7FnPNWh/9PZ/cax4/C0I4k/xJE6Oou+vV1W2ng2x2nq7j3Eemcq1I2OquBm6bv7C
39djh4pJe5nnbFolJ5W1LXGZmatEpp+swKOTwRGozlFzC5IIiomm3iDLReFoqbh2Drd7oXam+Sq3
l8DCnbAdV+q/dH2nKGTqhsjU6bWPTF+4XbVpg+yJzqNSbj0wsqR2EB5ENv4B9unmSAjWR5HXBDcn
JBkSJhhTQYcstRRQGJyDG5ahVkk8q7MmvsohOuEQd2SF0/WjJ6UkPD6W6ZIiSMfKtEBPDGIHJZRH
hw3Ic7lrQanncnmHjeLo7gQJehPz2d7TzU0wrM8Sma6iiCN50emQAZG4GlBY06GquHd8pvNih+WR
A41gvB5Lv+px9q/gqLvqPnf1WQ2GOU3s/LGdRUArTnoioeiHeks8AnCdqXmd+ruF8j/lcqkCP380
cgsyCBAQmZy9Vn3i2mPnbVYUKO15H1APJwOc2mrm+7cUP/Rile653JlrDaSq3sPrXgZzsk+6gfeh
+5LBk10NUTnGH3whVIrs/2DDyibAeHnpywP+DnmpEH00JpUJF8RllkdvHl0veoJr3jxlzCSoF72T
gYFNSDo5YYBsZS1JxK3rDl1t3x5HUHfeR1lLe8n6xqsP4h+lGiZHzliovEuY1H4OyJ1cjzoVjQsB
qOwrjmTr9Ls3RccCS+oymmfiLUrYzLNBEtGNkI03IiU2EczpOnGDWvOZItaUewKhSKHtk5vKESr2
4kKZ0tIFFJVqv5gQDxdleTvFoVgTOtHyxjBR1I2Nfn/kKDuB5vGlgOsyJxrU3ztxo7R5h9TRdwbz
lDL+nmlfaExHNzbrdYPNIg9lKmWvq56RZvW2yR+4P8rdfYGj7Y48NaC1h+QFoy/auRinGYSD8h+X
KFNgPTwn1e4hsRK+lA8mrtkH7gqJw0N1pgAlX4bdou7meU/WFz0I2uecyo3P+74pF1pYdxQZvDx0
VL4+xDld4A5Lg/9BtYoPdWsTiKmDGQSy8Sy/mLe3/fyPwNzqwstclXNSBM/8dfIOCQEkGXzkMeXw
l+yJlGmIv2A+rMxevm07pSWUnRZvtaOA7f1vtbbkcgPnLkAompdRf/X2ivoZ92YwWghrq8h4vVpx
Po0DWEnHv87m/EJf4DL9nZw71KVdfIV3pi5Vi3WMYjP33O2/oxAwKWvyz2DMqp6JYh8MhmqVoCJc
6qTZ2iZ4mxIVYj3x+Q0y7ygrPTGZOLT4O+HSU9IkaQTg5mbnsfwD/gYbiV2NHwY5kZM8n+ovDNJ2
IjtYUS+wSek9dTHb5tMjZB2vuTQBTlKtWgy6k2sLuQ68Lzt3wKp9DnNkBjivPrtl3eHHkpOIZlQs
ouBGQvzi76hQOz6vGxx5niSRTAiiM3fbquvPg6lUx3POchdfyJUvH80SYeJUq4Jx1zqZLoqTAfcN
cfNULHd0jIATP66Q/nfq6yZ7DQ/qvxgOtUV9ctuwm7H+Y7Z1yleUX0pqxrjOr0Yeba08DB9EPX5Z
oNqEvUh7EMxTSWyMmic/dfyZ8LP6r5aPa2X3/pYQOk+xpS3Xo/TD+wkOpb1UXKsuxh0RLSNhqdAE
oZJDVi/5COnqH1oDtV+nlq28+Q2Y1SHaefcCxlEyCj1l1S6G6tcw1LiTlhYIH6tNP1jjWInSMHlw
aXCRFhPOQIJvM7QFW/CLpB825vZmlRCl57rSyd2NNbb+JwStHmMjAoconfpqqvQkMgJOGnFng3J6
FWJ9I48l3ozQYVaam+uoedfQqAltJrDaEh1kub0Glem6JutkfjhOx/T3pW7jrO1OPSs5Oi6nwdJg
NXDLxg4NYDVOK0WW70rRvjputBke91XMXT24TVcuYVaqvLqSDNawrtgaiz7LhPtMw23zb/2kVjCg
gI1gTZqV7UB24KHsxEsM+xn/bBMMAoBFQyLi4PXTW/NWCEde7vhG6fQXvDDdvMc5JVIhENwv6HJK
n3JV/MLbUEjIc6XpVN2pLF7wYQImZm2ziOdmcjIQFjxBSbmP76A6iNBDyycHU/MALBfqLF9kfUjq
dsqvUTSgn4IiETBrKZj5WU10RhluYcoAM1+VEKf4/S9iBpe/zIt9wkdRwG/wr+BIAm0sH9+Q5wii
2JA+ht7HdONFrHbu5R6uIcrsmkh0W7Iuug25ZfRQanaP8vWl0eZsx2hImDFDC6B8G2aGvuvn+jec
cu4D48Pb5d9vj5qYKiD/PP4u1OesfEKmLlazFyVB4jJhTYu1BINJvDNgivwIyd3zs8wTO4I1iPj7
23yTNYVP+YGgoHBwZ9hszQcfwdix0nprM4sxfRmqVh7bCgih9LehqemaAfdN9/3/rysR5/GS6Xj9
WG2It+rRT+29gNOa1Rcxd+k7oi8TS/LsnvqT6ymsALH0coaTp4w9yrvg9h7wAMTjMKecs0pVpYtH
CCP6Y6y706VrM0uAHVxpH7Ej1kejMbVvkQ3sw7Wp99B+XSfLGx60amDKANFYdc9EH6UX2V6dR7TX
70O1h4vgx/7ZIAToG23NAoar2oUcK1f8E8XIH592jCXG3IuJUT7d9RDhFxjx2EMsyb7rCdo1Taer
eP3/2MGe+XRqw//56m29qj5TYsowWpoOL7dtir/Jp8mTuULeWdyOIXDd5RSsVahWNvK9f1nYQ9ql
oChMplMZYaIFeMBomt1hUcar5nV/Nm1fIcAnovii01NK+kc8A06mUe8z43N3eLZnXkH4JpDTfuzu
Glf/hMkZaJbxTBk47M8ArUHz+CuIpIKxw7Do1nWfIABqK2BaQHZu6FG9hcJ7sQhgp7txDgohq/M6
W4tDJzN1Q/W47DaYHMCvyHtbf12XSDRUATp6s5i0XnAYPnke9FmOo4BuYJ5HY9Swwjh/7RtC2xQO
4wqkZ9x3J/hXP4VjX9qvcjdWfoHYsIED+L9csQ+gWMujjdEkcaTC7Wk6JgcnVEQRKyN47eqnvo9Y
SsyrsWthTx+VJ/AMCgiRcv0X+Oiu+moKgEXcwg1866Dnse2ZHowIgGEmavPsmW/BQIMl2Q6wcCOD
EW8n5TGI5fRqhTycXSo62aAoh2O0CUg5OpxlMHuL+T/EjcNSJeUhvhlNgNXxwC//x47y/EMO88c2
Qewbx0YRu7i/wCiUW4JsSZTMLNXEh4aHIE680qgkqr54uyfH2dsufcgKIFkK7BEulq+eW7Dqm4H4
+61Iy2kbHs/JCP+QBhJ2cg405WigFNGaW4/0j0s7bglNGS3xWJ25/Uwn22j6baCBJuLjGgnS7JFj
Ybo/EMjF12EWceeTDCbXlfZsgJIuKvbqwkTpnV+P1EQMoKNUijj2ZpLHSV4bxdVN16ONGtA+7UJN
kATpb06dutzH7APvfL0XVngTU3kQKiXEVnCZJuqu93Dc7sqwDwiSOmYap3yEkRDZXvXf1/It6NK1
CEGDgYNex4RIr2Tuh6Tn6f+/DsMScIsHUUKvTOwJTzbZDValMQoFydKM44YSxhcjre3e+0YhSx0J
SakO+2VjA4Rxc0MwFelQujjfWw8ZqkB7CHjMTDDkN4E20LliLtfJXPEX4u6EW/mymfANYctsHD7Z
5WHe+HqZAr+0ZZ3fY4/wYb1L7685Exv+K0D0ZYZ4zR0Qg8W1MLhUi7xl2spsRMgYuhmQWToR+hSk
pTPGx6EWdPq259fx7cLXqpo/gr++JcU92w4HQK5EneJPPHWVPmMUFH1eos6EEep96L7H5N1XZCzN
rU4BeZEiFh5QNsKJapMIGs99DpVssahh00l5McFyYeZPFkUJTEy9JvsXxs/tFxr6qtNh8aEOpR32
W8KHLsNUHdQKRFbV4LKXMbbfm44qDUTPJQM1IdmvpxNDz0o4L9IKlBcYX4q0jHmMbSJcZVTFIGP9
dX+RB4opTLuPnWYoObkUkXnyGFEPQDEYQJ0kpTD6gDfZGHYaMtmLGNQt+IFWfl7HdWX5q0fJJ9/M
ysGFFeOjklgKrLafenVThwBJl2bD5LMSo4/1zi2V+DYNd451cEW6KTtNfjMZTliro6swr3JV/iEr
z6WcTXaRnBmC6I1qZNjpKuRMMsaLVmCQWbddcVyRGLGWQTaqVDiqc2I3ZykH5rbylRMEN9ScyHOn
vNxJe+COwYqj7tHYiWy1+AYX+wh2UQ/E33/0NoxSKwWgnl/YNOb1/xwKHcPQ/K9IPkPBKLeAiVPH
P2ufj1cSIaNJeu0dlUI25Q92ka3NE3ReMDRCRj/fKpyzZyeFQETPwoUu35ylZ+93GBiNzIDTjeGX
u2YxQZN16PqLsaJdc3aSs9b/2VcFPfznGojcNDFANidx/MAPCIxECleu2MrUkactkcrzRZ0ThUcR
V7XES6tYUtW1IXnVMW6y5eG0mjR7o04VVH0KIWATanuWD1OwG5/E0WFXinq2ycryP2XsdO7QC5s9
VSzZqu9Jphg5/DNpz/bDllAoffpxsWpoDw2NPeDlUCKZRp94UwVqinjK0tXOIV/LL/F/Yld7QRjh
mC41sKynmWCxFSe65C/J3zqEYyKhhkyf+xxdyDIz5+XDDYmA46fBxFBoTgdV0bMePqHFb7JdZNOf
MnuFxBzsPAQimY1cwGLDrUIHCpYW0XFKNoc4tcmBOzL/ozWgh4wF00Xg/ETktBJrZwwIVioSXiVi
AfBxbGL4nwmCg+ZoYE4l21N6ySZA/rmk1hfSStS1tEunSSwkfyhv1WSDVyLBo49xx6XJa4YnQude
N02pwZBQ2Xaw6F95aVioDLayISZ9VxnIVe7Q/PZFZmWYEQvboerdngiRF26g3RLlODBhdjQQzhmv
qQGwk0p7W0WE9hPZikiivOV1koVDUYVQGsWic44eajOGtw0uDWEZH4hY+t3LAJWl08YVdvdHtWRz
PJIC19yGRDkztqADWgriuVQp0F90MFZEdXa5KM884zV1U1QfvfxcP/WQfFX8a/fcBZO7pthVh/nY
eVLMm9HZl+eIAXnxzwxSj1hDzaSK8EI6tNSPRK3yWwTfSBbWoalDyhqI4TBcjFDsfMdpuFS9CAfv
4VmvYQdmnmxCoQPRaQRmMj6hl+1q2gt0BP9labIwjfdFwVEtQfY05T2TjHIyGJYt7PL0so0NB60R
p0St/TLvYp0tLMHQVmDuMsEv0VLs+zfBJc9LGcTQEw87AsmVGWoqc0t2FuVUxoD8zkFVY7fSMDOw
6qpJWxL4IPH3CX6fPmapzFjlHckNrDF399vqX0nT0T722rZAZk5W8FEMdgSFJsTHkmtus5nxSqQc
IZdJYZUk3rB4EwK4cDSJbJK74AftizFIrrV9xL0ks3LsY/5zDe4mN5pHuzY7VgV6c8rhQP+gQuH9
SNAaTYFrbBWcwMUY+9nGZPdIw1cd+AFP3zb5Qk0I5fueshBFh5A7kXBLb6I3regx6gXH/slKcABM
BCv9S2iwu1m5iaTvPbLstu2PyLMMEyv+c8xYLIrRMoOESQdWlwEmBiv4aYyiLwfM7Hmvsjz8WlJM
nMqWjy/ZCFjgr34I0ghwoG76kNsVVNLozcNJ9S+kiPITQ6UulsIovLjET2eK1RbQf+SWWSZ9dnS3
DfsiRpDUKNrJbm919CBGPuck29wrheoFtsL4Np1mHP5tiUTe7KVHK993EV0at935R72PnkVvGPgb
UEJq1rqQxSj70vxKXole8hINgPjM1VwO6h7sJOdcUS1y5ReLvvGe9Mg7/VxloVZOLe3SpU0bV4/b
jJanu3pebNcwKEGmSsIdqH1ZUKVoMr6ZfM5owIB4xW06m37heDM98DHKj/x8GgjIiHGkNA1ZuAoA
TXh+wSBpM8U94UTRPP5/hiHJ1N36cSGVH9WTo3DFMkCDj4mzTw3o7RP5dmeTm56WBUWQAE2B1N4a
q0V3fyIVo/BtAZ5JRugkCYpsygscirMR0R8Lmg06wPyWCRhSogJfmgvVkp1A3F3hYfvh46nCuA+O
iaulqGO0nKWZ+j9SDhl8/qX9eAyfnT/ieSItFPNPw7mWEO4AwJV/lcrEJzS4R0vbzFvaDGRMfavr
ZmUDs7j3rC/dNk1vVlv9qNgbi04OHpp8Ka6sATJphCaqrqdO47tRWTxggr0D6TVpwsd96xcJrk+q
Qkfd5pFpCdY+vndOSWT1Ly9NGrwSLq8odKpNtgb4iVEgVEUYPeFXBI5lH7gPb6hK3ZF9Q3KRH52Z
CxvB++S+COzBuRQDStQ9OU7hCPBUXNbTsd5O/EtBB0bOfBj3HDhGdjAmEuvUweNtvQh2IKmHfKFi
GRcWz3F4SqL8dVrXrJDinEWJAFwKEfMwIPlAU3DsIBKAxrOh3SB/p5RoewvwjMUiBj+82ZDUO1Ld
ZPX8K1Rrpd3fWVt8aZCTPeuDcm4l660VC1b1hUt7CUf5Wu7xSBPe4AG/lO0yZQcPaoxx+DD281Pu
1TvRPa7MOq1ujagVgsnnvCnsfgVz4P+q3UdxScEUfZ58wAvSXt+964NmKu/H4h3k4F50wHHBjYsZ
1fYX0bYYPUfdaFX8BTMO+Kbal3oe9a5DbSRCjHtGdzowpv7Qsc5Sj3f/i0PkWXQM5J4aXlgJcuXN
dp/4NheFFYAJayGpTAatmGCQjL8/iYxALmD2OG9iBwH0CX0+WIbQ+dp61y+ljbGC26q3FiEHE4sA
EhKdu+7tkrl6j8fwnjoKpumf/pX/a+ssOu8CPBoPYODvCj4Cdg+zOEkHX1vRlWTXUAxzgwy+lES7
HjHeOesbiHis+v4lkTEjGbfRlrf3HCZzok15dkbIpVPrMFelosgpo0dRiCToT+ZOh6DS1cge4zgi
T6FXeSX+JcbpOFyG3DdtsMPM0YQswkn+TA3ZRWsdbHgRCWZUtLRIKK4fGVxaBNJR5BDQNKU3dlgi
VrWZeSLAOiiK5Ws82904I1U94eegxN6qDaOWQ0Wwl/kC/qu7xVDfx+UvKybYl3KkBPagVdd3oEih
2EDHenoB/X6R6PstImiv/d+hm7FgLSxgwLTEIrelwhkZ6Y+M+9yJ/fV29YJcdmQ/eREScHsXmNt9
e9tzyOGAR9ro6gABQ9Ku8kexJk7JP7/uLsHaiBOzRTeNA2fVNgNlPytZx5x4lXzRgnxvXqfZ6kdu
nmJPt/HC00FgDVJZYLQg3OSXvOTFjAn2NkVxLVdQ3BdvRaYlSJhBt3lsjCGZeSPAOwM+W+rQhD0l
eIh1TxEfSxqp369GPWwj7U/mGQb23DkOo8q6eszBpcNkkvIeuLtqVlFB56nMDpQvDTIHmjU3S27q
MXKtFH5nIa8xHVSKtY7tGE1J0Ne0gFU73mTasdQ2LCTNVT6bFXIAPSU2+GvNY7W+6JwoFlWOvi1F
ml06uzui0JTWAj3ep5uPwlcbC8wiCQscJFLzQUWuLlKqjcDKQ4KWDyr9Mlhb8Ytyh/mXj/a8UjOP
/woDxJ5cjQtVniOQgJSO2SVbJv9WYDgFCPYQte25bgrC4CcfKmJcwCQu7FAt7IxBbeOuIpzOZYMr
WzZpSDjOy111cjAKloIsABIidrb/wW7Kc7UoLvXY0Du8ldawQeoBkf9/an1yHG7nYgU7MRHeg8E7
FBe11nz+zQAke07rfoXutDHFkTLAXz0D2Cfrf7l+A5s6RBcL4ZIHtgPSO/IO/tdMZNIqPSaqZJ1G
CLEKjAOPp+tjTijGurP4KQ7JMpT13GUL/XBchj2HrwbMuo368Gh7GThGJPxL7tX+ko05C0uTQbMy
tdgLhvWaTmSlZqv1Sj3kYWTB4VMJ8Mr+Og184qhES5KDDZaT3tiuMK9kf8HEB8lcVgrKcVTuH/NZ
Ztno0nuESy8uVrqkQWSgaNWl++yc1wKG7JN49pSzWQqAnFPxv+jjaZYBYxfkbXy5cHZmNYwxhoWd
2RU85tnJ4qb4Cgwo7RAf1csYjBWN9BRa4TzIO7W6PP71bTHGd81Kuz6apIUDj7ZJt6MegVdMlvuB
DhjWqQ8XzXkeomYR8HVU7b5yaSc+AKwCGUCzI1uG7yRjNzjIqOArqFw9FvfgDdyIgDTeKYQOTQDm
6Xuf8vTN8x8OUgrzRqUuamnC8wVx573ITi43hDYvjs2DC1yODfmpt+CsbyVw5xJFGjswlSyllALo
vxMNNewQexcbs/CwYIJi3GyWPfcQdGzHDR/XPe6udONsziocHWuiehmmKsfzZPf+C5o16LwWpBrL
yVmILJFWAv84OY/CIeC+xWeblYB6WSaiwqkIpmpS7JuyVoqP2jRApEjJQ6Eu/ZLUHCQfNUx4ACGR
ZE2op92e/8aDkmlPmKWMVrhd4Fj8fnGmzRQSCz7GDMExnVPV4unNGebRCljhQMPqXLTon0TeLtAK
nttI6YfQkIq0vyq9IGH08G2eb/8U/KwPa8SYdAjZP1gMX6FlmeWUvn3Bf/kB43pPpT0HTw6xcWvK
Dz6NeIBBm/1a0joZVW2Wac+jMW3GQlIJKLawyIk3BkF/QSAFed9B5sVtcfugVQf0P76YyoiUz4Sa
tCxNYRUvgur/PbLVNYtoWS6XEKAuoN4T/E36jmaTujVPZdyor5KlJyd13070YRpBfXr+5y1GTZJH
TFdFN6ooych70TmL4qSY7b4+fSadhtjNdBIs6SX2olJbIddq4dzJjSCICoQp4xpgrlRpVdHfD16Y
3rfmfLBY46DwqaGxjyHqfUKYOCUO3W0dOlW9qg9+wKUJ4GHGoBNsT7HbYVXmnyKGSNuQwksUNmsT
vO8f2uGmT6hmyeaYUAYeiVtHMT1Oqq8AXra+04fNZaTTSvg90WSKjepxZ1yonLvGnTqni2IO2T+c
ty3f3/d3mFOSoUoCPde7r669ereHgO6Q6MIwNJjLYi0eP+DJ07bKp0C2m8i7E2iFMRuvD6SNwU0I
ylQuU7wxqCD1oOCpz+57SMBoCGJeeGiRGW1COgEUBj4mXRoVaTPGtIgDV0cSEFeX0R+3vga92M5j
EVhOIygKxkCi6kgNSlNGFN9RXMEDXB40L/3DJ+Sz226aoarcYKoXy+g0pqv9Kghih/xNqEXNYt97
4fdfdheTlX5sDRgjT2/8a2kZc1pMVhEAHs4iCy/ar6HwMqij8N/nhZlUlAqSllAd36VEx5AaYqqt
brMPIqjnZmIhFeBRRMBQbld9hPya5EKR2BXF6Gh2IJmHZwlrQ7vfFXrxVdJV2dHc/ECSK76+8VCd
7o7pig7Lcwj3ps7DnIUlS5XxU20gGBej23vdrwo+j1QbH16Yc5uQZGQmJtZhWsWmQVHkl+fYMRXm
uigzW72rDKTeV4w0x/Vy8aMqPw+LpcXLmdLXdJgbKIG3p4YmxZvMP3Ml0wIVmNtIXXjVrcrNpG0y
emw2LVwd1RyZ/cx8jHC1j0IuB5TcW5ZRipLm8YOnb8PEWDxRNJBIDShUKilbW0pz/XkERcr4Q2iY
VWQC6II1Gf9teIfi893SHPD1rE/IjOjRVq0Ews8WO26/+UJE7Hw0vTZ69nDALe5BuK9HNWcVjAXV
HgTGrMPLgStfjZHe8Eip191fcD6NavIGW7dccTpKxag/c1iBCURc+/gau5GXJP0vJ9Yrs4Kh405O
P+ynxA8Ng7+pHTrGi1r8zHQ3nocshGMrJxsbrMLdG/DCQIrnfweDXKbvrilWxfDVMZzisMu0YQBz
koGa1A6TpV0CA6DxvUYBhnY8ncL4ey6VmMDi3Pv2Eg/GlgSAHrAbcaTn5yzHGP87SMvVjYX35F1B
/FP6LoSAGhxJRmP05794J665tpYFEUUjd2XrWtQpy7yVC56UnXh+MU8PbCYYmIkoxt73EsRhsKyx
Rp09yGoUQ6LLgfGLWhYQKcb7TERIQH8HosW0DWRdKNEa8anS8FPh6xkw8TQLp3XJ0Ex2UWJe9Ksh
iULD5NAP5lF9SAEfx2oKNCsufhYPkXxd60gIGKG0j9Om6720paNPnGPDPQFHNAyk1olXH4HSBIM0
PJXngwfRGYS7/ePHJArNoo7cSR+p7Uveqc7Qzt1OfwPyBj1VTkWXr9L6l8anWeKq7Nu2tgHWctHZ
0zK8RjGSJjz9Pt4E6Ep13d7dMxlt5zW/aBCrujWtZNtwFMPzoYrRc6uybIsTcHUkuydllsSIc1BJ
kxoblcEMHBXd3K2W6e79XMejWS0fsGtxS8hMsnjYLfVFKjfU5S10Cn4knOTYHazlIBD9Z592/ebW
JgbIGIUOCLUHvuf8I7f2GKmhYkekYBZ504b+sM7hND42YRHXJDHpZsqLni+oZnz3PCMqPHQp9pfM
n6+nzHL1cRQwmC5rhq300LXZiCPhXCRbUJW6NGbSnfuic+e2UT71hxDccMuJtc+0vsCiUY2GvITy
8CVXwmRTUtYkFN/0QgXGTwTSVrb3wmMnvWMaUdo54qBwmZA5QEoe7PieRg5wapFRzYv0fSy+4rBA
AqkH9XKLhH/Xq2qxMpUmYUMsTI5pVLgiI2mGhXlbQ/H2M3KjyfJrZINNXjTWUFnMHfSqjR6/UPyY
HBL1x6kQQu5vU8+DrYjfWU+E02MeulXArCZigIi3lCU4mkyyHVSnqer9IWStjB8FDnTy0wZoC32l
8stPi9XEEKRy2Ghf2pSgJ4A7PTTHoqlhDhP25zNYb2ZYfT6s3fdf+4CMhPRWVIecVpV+an9vULP8
17wfu+BGKXcTaHC58pRCOLmC/+7IVotIK48I4sD+uA3ByVN4J+MijKRzO2slpiY2tKrUE8hhRkaN
98jow1m1Jy4Y+AMlIPPsZOrZ0QZcNeWxnAnFsBYI9JsjhuRpXzLxr46jzsmwXgqkaoOrdNwDNP0p
PptMfsxuzW+uqh1q62VzKqnyK0OYbBgeNBoyd8UmgxCb8VxQoybJ/wOpNo8FIJYK/MsZMKpBo6c4
lPSb4f9TxmpaZEV7oI+r1I0f8JXy7ixU0hyDBWQkUM4oxCXF6M3Zj6V9iP4qM0H6zrWCC78YtQwZ
HA8pA9ofkcnoeDbWSQhWT1wDoY/gkLRqE3LMNYHULjmGDRcuub0AVGC7NenXPgIf8/qCOCkEZ2QJ
w2azeIPPljl6vU04xki/Dlc/yjTNFtT42ffr42y5Y/WF6JUF2PNIBqbYYD2CvIwHBw0//hUZOZ3g
5EwCo8kfbRIe9hHAyaw+Z9hRfQ7Ay4LG8HTo66SlQDy3SQOYu8pkdmA5MDxB3lNwSEXdkjMi8DEO
4QEs6VEeyj6l3OudI2dlaHqUz+dEhoj/ak7nrk73JpEa4IaeXoQ4Gn4pey7OUFGqS32zSkhx6m7c
AIFwTV+4Wwl/WIYFUUTXmtcswNzn3+mJcJjDQMhrecEMDwbB1hCQ/uE3cBSYdeRICTLvLyJgizAO
f38EWY3CS4HaOBgyFJvyaDDNRBwXCp0hKdd/nKuiP8qD1aV+HBW99WCV1AL7KCeieZewSY6CqFkz
D4GHZ+TAFFWI77QtW8zh11SEk39eXSSuQiWHI2BVvUuIaakRH3catUdM2t+ZTv/Ou6n03qVlVcjL
VixfS6qAdo88PAhjAIWM5FuUduK5Gxz0PBKF+pNWBuLY3bA0/a83MEqeCIPXCm+ZQY/IElKqvZyW
4bSWk1hQvKixrab5Ly38wbT6uRdIx0D2lOZs+6iTraJ6lAS7lrGT6AUJRwIbQNg3cUjSboY+t5tC
/r8lgvElguB0uH/d6oeBgzSihcw5GCeF8zhRfaaB6sSea1xC2uko4XUcux5R/cEqpC7l2CDds6Ki
v1xoShAmnrBZVH6fW0an4K43bUeK7k2b73KSbCPpVn1b6nVNZVX+AvJnJp7dXb4m2hxgP28Jh4gz
7oI3PG7hMS53Svg2YWRyqdXT0bsV8O/MgmmAM7Wa4V/wh5R3CQ2/t1dWgpDzBrk/72PEP8Bbvpfm
8p8QuTqMi0TJyQRi2wMckJK6UN1naB4paEgzHOwvSbGMtz0jlwuTFuo4NDcu2bxcM24xpao2jKwp
DXaRjg4hSlSlJzO4i8CqToXDqyAgb0J1KSUuGxjU9TLcv9T1o1+MKv+L2DyslrDbOVEoKL0kay5L
YtEiv0Pz/XfXycJs1rtnksM+SrCE/GzGGDS47zt7HK8VFae5YsnUNEFjDXvN1zcHivluRItH3bp2
GJvM8r17jDZcNYV1qm0/8T/MnAgXBAvT97twUuf5GT9eD3Jv8FOZg77uPx8ajbkm8c+IzMuqxNKj
sDOeO9eEQJNDmFlNrf+pHBnCfUo52RBycco6fVCuNRQ6cDbi5QsIVssk1O39Sfmg/k4nYPXMFwLV
B5DHy4OEMz3casyReCzKIhlzqUCklmUuLy1WMjCm97oNNupOMSLfdheocPdjW2P+4D+urzc9erxn
3gAUYaAkVJHTtD+P2MEDb2LZgYWy418Pxhp3hEBqInoX7m0A2HDUrzlvNMsS7RDAvNFR+8cSUzP6
O/s//rDspcqO3lQY9nRjW/2gHRhedffGoM/Qa+PYFbyysNk62MclUZP7aV3UocwQ0SW4r5go9+vi
fWxbFGu4aroAMVaKu9ukZfyogll3+FD6tJj+Vrl48LfVit6OyWAz2vICwl1tRDw8gCuS0kMGLVUX
E3TsmLpB4s3rzpsf0BfJ4spQ82JsAQ2Vq4YnY9Bt4jx2uPvQhE5YpSwp8ucBJGZQDEdm5Y5MjZgR
/4aAARRMFHVETMlyH/8F5IUJe00Mv40dIoodJn1bxbWOzh6UsgG4zCWR7rrPuJWaSz7LCO4lvOh/
b6/aiSDOJAaGHD/YlTMqNghNSOV1jXW/gyeQ0FssRBXMI7FB7UygVWcD0MS04JcyiQwKP5VpdDmy
mfXLiJhge2ALPjkPQP3aXJbM/oGA6kkqbpIaDMLd5bz+YH+A2cXqJLOqSOzriilml/EGwIB9tEZU
9nMa6UPZhTUHeJzOXBrPde91hq9B2U3L9zGE8t4Np2NBSLGzTOlrjVP8ay0qV93UaaqsaqOQH4rf
KsC55YYuRZd4xqKXZGKW8csLBZOMUI/AGXz5/5ib1cgOR5iipoJiPTGopuFn3khjHH6Dm7PpyuK4
D0nrDX9ZsQMnbg4z9c0dImxWK+HAuEG0c9SelZkio1371Xei+nlVxretBhsx+3FnM30QJOVayVag
HkOe50VwuRhAzCdzwhcM2xgw9wk3EWX2sjBKuDa3TvgAZzs7Ql4816lEVFJyz3SDwrqSAkZRLpFB
1CBNccBUP4P26MNPa2nXHlqTXlO/yB/ZUjT2oKXsY7wNINUk9vDwil82z+OsiWQWJp+sFCNIyIbz
m9lnzRKI6pIi2szTMeGZIpismj/gnKRQ9/A4wlNoI3fy5BekiOWveoC/GUESqT/YOp1XydDrF94p
F7WTLmQ9M9dccGZyugGZwCcmszYynjqBH+HoSdZ3u28nLaBqicxQNvJhArH/xroQ0nuGRJtF3Iwu
5RKPbKd+IEQ8WQxGuR7aaN4PvaahwYIb7aOPXetjxVwj/veCB4mlFjsSVptlMGSBRiBYQ42YJuKh
6d3WyIWYTbuuouPK5qygVXu6oV8i8Kao/vEGFuwzYjYpdiZmbPParSRQcLd/QCPfcZ1xYGP3PbKG
ZP7VRwOUzcg0lnvnSvCOnH459UCOswEDY/FEtyuFXpVPXcGXvQ1eh6kpyOMDBRe1ssoPl754Ku8G
FDFX5XgExdf6Nn0fF55r4ZxyTIT2luLjCBO8nNLWTJ5OvBt8em2YFd5EmNPJkyP8ftCOQakSbtaS
tuZK/XX4+Ao/oQxGHQMzKlzroyS1DJlXN1Fzdr5I/dxPaOc5tYGcUnp56hYW67mzVBTQ47f+t/M2
o6C35xs0BZ0dDgb4UAiIfr1lVfQSf27YeQRNna0usfX811dDQQ6a3pKXCPpf5im7xxmFtEwu0zYS
bTt5hqLomKyxXzNXBU8HEgxq05//xzdFg4xvbNnDig0u35S6WfWQEyLEDx+sW9M/f3gBzaN8y95R
Wwpid/aXN1FK0pfR9OwnKwOfFbkzz6CiEeRaEmA1JGtSfxZUovW/w6HYsdgvjlHVd7ehePmaxXZ7
TW7Y3yMde0GynrqFhYcDHN+GvtfWyBug/KZlW0xi/G6cCqcfZQwQ2gqjTO85iK7ZJJ7XjHDonn3U
kSmbPR/SqThP82jLU1QonnqjGLLYEtmcw87VRW3cWIPdjjlK1bXlAi8FQ67OGRxt/wDy4nmhBZlJ
XpL4pGQEJ3F11/j/ZqsbMFbDWIIyH9HChtYxYAtsnud7FglXZLjhtXbC7PJRxT2m9SIQ21Ik4mm+
y/I3/WkSN2xsnMRYnS/b6D5fNQBFYLmvGGKJIf3Up3hDw5kRFtfqc0V+B4dKRuY3NlhnV6tXOAI1
y0ZRUhQtQsyepGic8PtSEaMTKq355LCU2CJ93AJj9cJH4i2VSoBA+pJDTt0i5HFOSsO9nJX2O7vf
REL0TI9McIgwEdl2y+Y0TfvZ82VERIZtxsPDXP0LKesDTWv8rOqVtW6Ujsj6LuHFnRBM1D5UEJ3i
dWqTnvx37SNaD1An5r4tdn1fCSsIXvJguwRhtAGfzy/k11OqSPUu6xkloZZi/tZaM5/KubHWEXma
Uia1r0QuMOC6dDqLgknWOC6IlvzEfN4cpX++2BH/Sdf4Vow4/LOOqv/ueF9L7sz3/AmsukXDvfRb
wj8L/0GOmc9bmeT6ob/VcHl5aLkvZuIE8MZifXMRo2KXJ7cdYuuYHXEzi9rg+L6JE+ChsbeEMJ5l
7/vELjh+Nq6/imLIjP6GHbyoKnfIIDkvgvOsFKCKWJ7o6MhcO4uqw0/AR8GaWZiKg+cMHRWAVOJq
ojwrJzrYH/0/VgU30vqb1sJzByOjTlClo/KWJ3izjMbmk6+BXLIZ1ekFNwmx792t9vsCvCTqHSZL
yXJWW0dvKUg9Hx2VDP9qwXlnk6OLi3H1zgeU8Oa7eBQxawmwSbGFcz4kje4S1c3tT9fzb/2JsI/c
lap4vgXC39OE7cKEx6iEDsaGbMbV3zxqNoYJM49QdOXevYfjGsL0qh5TRo5YXe8ZEkdcSfUvw+wm
l4waYKltjFZ69aGejJGQBIj+gSqNmiVpEx5A/2dDwGTL+qiPOxyvRjjhsUBq1yBkYS3UsUl20g0P
h/5e262OPT7TOXr4mrMiJVisxcRx/6gdxbbtfqiwo4weBLauC/I5xgkshqDla5FVL9G2BZzRZ8UQ
5hu7Rv5VBgqXskNXsxESzcjShOQj1JazMsco0xbbl3VvaypHj34M4B6DXYq9lIJ5QmB8KCIEv8g9
NBdAVcHBzhnL80GhBHfp5rGGrP0Pb6O4TMonBvy8yADuDajfdeaLPjfUmLlcPFUTOHk3mkAiVr5Z
/NhTi/BWbteVwhb/aVrJpQSlKrb0WUeda4EPYGokWUbikYq9C6zveqr4hLkaXvtzyKUSQwcze+hx
rSSMMeWcghDecofJK195WcAL4uHRtpm7h8OLyGq5RsVmwVA3FxJN+XJZqC5Y3sloBHzSoD0lE22S
0vtBE4V/cmQPJqpoBEPVxbiUfV0f5wNdGg8SImCubjz+VOdghvH3yhP/JhCzJRf01Brunvdxg0Vs
1+yyXbic+PUX31c9HxMVQe2alXIYuzyrDfM/XP+5ptav3Qo0gADF5LxbpAZy57afHShSQTZBxDzz
T7nmVRc/kdJkMrsqxAlH4E8mj2CBCZw+a/sBVpvEB3J2ACwflbAFx2fi2GbxyEetOt6w0lvQKjzW
ZfIEsXpRWrAU1SZzYATNBGjLM/DxirNOpyZXQD0SkBEUHVJ0DQivPVFIWy+zh2YNOxTzmwMKqPuh
kp4M3zDyVX+9wbKiUjiG+tJ+zI0qlKBqbBHOe9stMvV8waBe7DpgMwoxNT5r8KO86MM5ORE/foCZ
b2vilL5Rx8tSDgrmTlaDdwAdq63ViEpSVzTOCKVf4pcRsi4e1mtW54Zcwmnqs3sP9BFLKuSpkZC5
nHeBZDRquytglFFsJMLlufZQEQD+82CwWJRZfC1qnPKX53utk4sUlTwyG8yFkgFqfjQIVn7m6+zm
OVo/p3nXSDr8093S22k5QaMUcst1YW4rXVoFWAyycFGbYM5TZnlLbf3mUaeWySqvYlZZ4E1KGcpp
wRI/3soEbGcc2e/7q8dNFORfw15zWbQX7hN4Zj1sxYum4UEAC01r1YnBghSfyBvrAQAZxGUlc8Wy
+yvob+JK4KntUnoOLT25Ts9QjEH5QuzMhQljuwsMHFMzXl5s1+vLnDqSnXw8i+D1500bAocLkwuA
2l2pucoGnRKHXg6NFQ18jB+2t6uIk2A2Qf7Al6eHNriS3x07XCX6ViECxUshzHuenPngZhovB7B8
aszenO6XPU1GfmAer1fKKFifY1FxummkrQSWy4wV5A/DmJH9E2lnzLC/bGkTx/x4JWP4ipcJESiZ
nALuDfyB27hL//Ujy3LmPsvgzsx90EyMHXvPO0zQ+19mt1HE3X6s+oYBRw5ldy0D6q4LqjPtj3Sm
37/Fdq2eG4GouFAvXKK2qIG5Et8UxHla7fjMXQNajDj61F6VIi+ogmCHD+2wj9sJZ/MtFYhc3zSV
X+CIlI0XDQh4HM88VpzVZHGr+cZtqGSPO5GctEW0mTgJo5MOylRYJ/zX2WnmFP2Bh0dt+Vd7Vq0J
sgtCqw7kDMUTsQh8CLx6lMFB634F07nur0e1WlqcsrOSffOCkxNx80BRkU9awHL/KEFjLoV+dPiJ
1eKh0I/iIL2/QlNzGtwYQsA6mK3fwFva/sA83djXRrp2nZ0HAeZAPr4kG7pt3E2i/Q+9o/ng/0j9
HGUflrOegjXofmGba+bgIsn3rArFmsny+Nu31ZtJt3VUotJzCexI44dgNvkCE9aJ1E1zlukyA3n7
+Qiq8DbYFxijcWldniu+Q928E4L2FDloGTBzypqY3S9lv/Xh4U19wuU+bqn7cHumrCGvVBD5ms8R
y/u/9zXYET3l2lfX0UlamaN/KX21ajtmi9cmV18mTCJ70M91k3DcROWhnBcZu+O8C4t4XF+I16+w
Pyyr3r2RFHKnE0hIavOISPmtVY8KAVEqgiT19+z6wmRI5cRwPALhAC0g+gj2Q5ooDvIAonI6eSkn
vz+UCbx86qIREEuFLxSB4DzFksDHQwbTODSsbG79ahsVwQyVI9ZxRB878netWrPXs+iXkFP6huqX
0/l8Y9+UrTl6Ue0UCOWFINDYVmIPxHY448lC4hbKgYAbKy9J4ZW3tUcIlyfGUVpQpCnbM59Zz2iG
mqj06ZwLcg57fQzcrEDqyFwcvgd3taEXsnGe3IJPS8NvupQJ9y1oI4JzMSrH3JJ/lXQoUnVq4LcB
Qa5T3kUa/F10Eax6VFIg5zQ+XdP1f/g9h24SZmEAf+389qI+RLZLqKiAArFlNZ/g8OZmW+MusyL8
+jkx4/fVT3On8bqzia8+iuOaGAu+rKXuyimLy2nHyXj8VAIEdfLuzxInpsesL0Vcha7KP8QRMTFc
o1WcdIDUjGlXiKU/s0EWwSGiSp5p41NzZh0aorFkOR3pN651xsyVkiqgiUeOTHwPXgu6VcX5shAD
OCUghpHL5+IEfxNbrClUfr4XIM15qvR55mGD8qLLRT5jVAulJPuMCNLMMKbmD7rgZneH095Lcjrd
MGo1lWNW/RvFTPeXBIzgqzgUm0DZpoKTRFw/+pcJ8ScMvIpN6kzq4ZPfjFeCBKbqBLSf0/oOldMw
vNgzJE3en++AC31z9YUQA47HSmHgcJNnW2akPkkO87OoXEYHeFRKMu/aJ1Nw18G2I6K4qfBT2drP
GnjEAtVeOAYapfXvlTVliqeAm2u5K0GRbXDz4eoZ9Vxx6jW9d9MiMjUS88ZSbj63GWaiklxZxX3P
cCwjyk1yU7abAG4mEqSSZJAVUHnaNE2yxgFS3+lGVdCHeLGwtklox+Tys4u1Uvmd5hhFBKTLgvvU
8YmIJCQ2YTBoRhH+MK+v2Pi/4jUnPcvt8pK/7q44aYEAMqBL/2Vqyqg/iPOb6HOro1iCu4TmQxFf
uG2WDztYAuPo36T3jvLNnI/Xp9ldy7drUSGkUiCXgU6YCeQpAf16iD77ee8jYEecLdryICSGGhIk
XJr+bNRqKg2NYu5JHLDqlEBz++Fn+2gBIUYsTmUdogGg9/r3x5789vln5JhDOJJ81x0dzUeng6R/
iiHaGBfGBogy1r0ec9WgA4Ug67b1hUaItSkkdzTEdXE0FY5UZOaOd3pRU8T6pGIs4i+d1USJ7i0I
sd8cy9hNdxJjLK/jmYbQozFjH6ZtALGChSLYZvdXBR+JQDLEKvcwZX4/P2W9KW+gGTsqZr2eeqz/
kzvMGswe+IcOr/Rs2Ye/Z1vz3zcEPWJHJpttjidx5GOuSsXfL9JUodwvt7ZkTT1Lz7iKl4k7B22m
j0vAeshWw4v9wQvBbOeBxSrvloU2n4YJIvp42j0y8g0GAi01K3CsvOQSCv67xQl3qiBTqiCtt2nf
a2gy3nmh1RkPaSvMvaKUXsOBJcndHEnt+EaM7U6HqaIAkn5uua/UHVlv5oSwkbhkWdWCf4u9RqBR
128uXrMnNz8UrXJWZ9ZU73FZfyjym4uTj0t+7Uw/gMiJGfgNJha+bpNumsfGxIaucD8DXnCzZNMq
+XHWjp9UoNy53VHZY7SYb6TQusS4H9w8+5t1pJDsbt5JMrD6037x3xcTApe6y0IUKlvpRoiKLHe5
6/ZSGfQU/jgwdOv7j1LEAxyB64EkOjQnJu8hnsAfDWcPXoUIcOTN49OAFMrVxjpzYObkaKi+PPec
FDn8ygdHvJ9Mtm8FO+Tw1ZTkSyXRT6P4LmZhy8MooHSYt7qJogzOPKuVfNO9v2LOCnBWs6bqtIda
BEbhJLrNP5d1/Cpd7lztPriLe/cvGrOlD4uqC97Skb7qEzwHPLp1lDIVpEB1/wwmbvT+iYiXYJ3P
+52F4LhQxKbDIySBeLTwJZ4N+KuJr4Isq7TXbC/XLxwYNT+wO/a2gl61DK+EIeCLgWlEWRkM9rt4
dW85viMy0ChH4xZTMTRRyafOZbOwqMzmdkho/PrB2R8oyJitvN7szLP1dSHqLJ+brbzdAm0bGB3O
i3lF+lXzvMmSuQTW4WY38bt7VF3ssvTesMKzDl7GW8Wl6iisHhC+uTTv5WzMJEJooKtTJ0Fm6sSH
hn6l8HgVqzTq/iB1AVcQ6XqUt/6sNsag1GYtm1ls497xTIn7iF5y8FrRrcqaoVm/5ViuQfR7FRK1
BK6tTpODaEx0Yx/jaR1DUHrzadEh0CAx1jM7W9KkMJcBT5GUunuzxf508vrrGmoCDgjR0ZLhhq6v
ZR55rCFCCnZ7kuAUDatDv0KoH6CEFBlI62gyHPrcRodlFUz2Eif/KqkNiGGUy/HSUbMI3yE+a4BR
CupmCLRBhZ6NbuzbHA3BoBpKtqfg0lS96NL1q63KyxSqqJZbvOq6Xn5KAL/8uJwVUr8QxP9LaNro
WUmh/SU1zU6swW9g/BX+nEtuLVnlt6ys599k2ZgOirPu6HdxcGcyvOhrlnj2VUab9A78pRMxS8WH
icU/n3R5XrWZzOqDVMlXu2v5aOrffW3ZztEFRcZpJ2kpVuLC4Yl560/nA6In45lWP4UjKc04tbwc
WVWqlB0mzamiSrgt/lo8ymeXOF4Fv3dMY3pCiK0M+261p3rv8J7/Oyz5ySzCmaAzWqGoihJF8OPy
VSYPDyV2ETO9YqV9qNXb0/vQumWfKVRre8J0zT4KP8jzWnCBpRZLllIvwYZqBLoCeE0J3wLKWLhV
NyQpz/G8rI8Ksn3OBIRQLmZTkLjcEhMXgmlH6bio1v2phvJDBDJCHIiSAJ0rQ4Kw9QjB3n2bCQyv
gFxjcb2BmjY32+HBmIAFdg+vBVuGb/cwK/J0d+kTLZckQ5kqBono7dr0k1UH21jcMXVNHuOdVajL
oSyk3kqMwV5Nt70ybWZXlbKbKncEwMPashRtg28EfJqR4Vc/1CVtRgALMeWFmAoe+Un8M7ngoxZE
ya4PSiUdYu3W8S1ANUjI0lN8kTRgO5HRMoN7scUTsrXIVDyQkuoEA/3d3L8crO0R/6f3IGBzLhcF
jO9G1yUpttKclttZbppoaZ8jEJMIrDbHksbTpGcf1yfe3NxYfuxp2bXyyi/qZd9M8vi24FAyPR54
Q84v0w7K9NEL/p/sImYo9QOjuaIdtaUZjhtDy/tnIomBAk9Cq3KrqXSxP/v80TAq0qlbRgUz0PyJ
2EjECR5yR9GV68IIDpNrxUV7QlBsx6PSVTaw6YVndkLyvoTXkuC3vDpMzntPS2hleX+ax3+TwGyb
h3aNJsIMsKL/dKt3aG5UuKc52REWKSu8tU9I1rXuz/Td7SCQCltGT15haXrMqNklignr8eST14ki
lvDThNQhgD2XQnBC/i40cIdJ3RoIrV1UaqAZZdrvDjdHunh5cYWxjWsx4uOollHDWkRTBdRxC2F/
+xGjLwaaLyY+BOYvYGdCmxazxMi9QAjzV2bt/GgrjVSwxA0s0089RO2aaf39kv5/9JZKRdMEYc6X
b3cAXQkW30OAH5X7sWnxCxTL/POod+EP0ifL1zPE3W7P4H59hXmMX3j+QVIoa35hnvaAO4gj6e52
s830TsSkkfxHRDbG9xPit2mOI+a3UyvfodSJv2AL6abJntit21Q0Q7nhlQYpLRaLwYyWPXU4hagJ
fIOTt0/uVplTK1rMDoQTVS8q3fgjIjXuUTL6knO78tIYxCttjcFENDjd2Z9k9vL2UE6PPW6+UNxC
VewZ7E78nuzKfn1XERKdBwkh01Fa7sB1oy1FijZ5HPJLGhLQyAFojhTFeAFuY9LX6nlNSmJUjU3Q
AWaXe0N58WZ9Gz8NtAScaagQtIPdyu0dylwxm3MlyQpvljurA02umunj1Eoe5iT3Tw662qOl1s32
5QZSdZavXFrEZ+xa18CfMRQy8q7fmfTWC26zmPRFNsNLk8bcJLAptNpytvDmfia1wPtq5SD5SeBg
8uP2z8Y2jbjBP6Q4TJHQpOWTIeS6EcGO3AMDrG6bI3+Q1Am+dNvZp7+wJFrDqPZOe+aZ4pAImYea
r6QdQHdnDK8GBu+LLgwIsmcpapOh+SS+0ueXvtQh6tT6CaB6nSdCKA4iclolyD84f/jtpRA73Dot
Z6DjujDxlFYgUz0VatBMVd1ibdnocKYV6xUD9FR8NoNYSX8yvAWn2duU1ovrvurBrnHMxN51hylv
Lz1kdD/6nx8dwVE28zPMEgy/EBqD+qG2KuXsi6JbkpBQ/OKPBK8mnZr3B8YFXQvG7EIDvgx1UmwH
h/oKnIQJDmtuzu2PkP/cnoz0ugreqz6Ac7OPm8Tu1thU+hKVAFYkVVI1cqxkUxtKPOZvXrEiMoZ3
++vcoHN88pB8ZPxtErDnfqWtTfoXLgUdBHNZVT9srRpPVjrYFTdiOPxahRBgGxYuRocgYYd1m6Ca
FGl8M6vnspAP9Vf0Z4yCYo9ofz8Z0jLwZfkVFNBVAK2vCE5NaYKb7DwtbL0QStMYTgoHnRbQp+Cz
UZhPhmLp+PAPPw5Wd2aSpFQR+ZeXKlSNO6pNirvpql/iPjIyGFrVsKfTKzxLzMRz1Mw9ccL+id3j
L3bpj4UTMkO1Fus8G009Y+YSngjKthM2qa8gtw5LRliHcVpo9weLNdMLNNN366mNgZiY5knmGFSQ
4XwVDJBfUALt2VtIh7tUubSihVRTBSjeefyDV/khaH/wMM2Zvalh2m2uPNuPLbRlBTgQ/k4vaUNH
cxbqG5pTLXp5OtVo+flRmh6Ul+UVy1duqhsV/Vz2E+2rwIecJ9oZnv8If7SNnEsaK0hsVC/Kqkd0
pAaz6sV0uSoBUicsZJbj6hGvLTqoXu4/T5Ekvbg0ehVZDy8pkPGXyXR/R+03ZuqkBeVoBiVjljwj
iTWXBAupeCWLbc7b5JQVFl/9IkCrq6y7+8dIfJ4+l/QsXdiz7bUit4Jb2ehvoqaKBAWdR3lOZKkQ
m+Sp1IU+LRnGT48Bd5OzvvvawL81/dJj3bFrszHYEo5hAfVQZuyOX6Hu8iUqC6sKa6uaB39pC92+
1sFafFBlRGP84XOAdZ6ICAOef5LS4XlyorIQIl8IZm/IFOfcAGMtdYM8VN8e6P4fSQzS4it3gTHg
BIO7MZav9PCznnfx++oKm4NtxQmiana4uOh1Aig4DHd0J/tGY7gzhbvtXJChMk3LVfO9SO6gimwv
oycsm94EzDElCLf5Bny38sKqP6oycnIfvRglpOFDP7Kr23L9nODC6/M0WDz6YLPzqRO7yGDZ9L9p
6tIdXyvkR1/RKElyNizWXV6OyBURL9gam5aWOyTqUHxcdLphCyrF7/XH34SE90g3KK34KJJmXt5D
seYXn6L+FjTdYcTR/P4ClbYNNpaXM8u3KUEsnwbJUrCFDsyTWPjEUwoer4u1scCskRnSnDxfTyaG
4we8ftjKpai9+WkydMDtmdGln6swgACqZk+7RzijmE90YbZHyhVUIO52zvXkTpvsz2MPtIo150Ak
5PDfNyK2bh0ZwuHix7fy1N+57VDJ0FHi2jQiXV8jprygIypGcOM6pGkAfH7ypwSwbDKYYYT71kml
s6uaRj2Z+H7W3vm1VIHbKko/HsBegvIjjXl9V7aN1OqTbGYEG0KexsOL9cE8M8QhpNsxHmNfzhKO
dUAs3mN9lm9O6Lt9pHIzWrRCe9uochUBAxazaT2nC3+BrmgSLxAUSOfysDCZ061JSa+QoS+9IfAF
pVsiexVjRrJbdrX3GXaxlrMBz7llROIb3bhNKw8u06SKVb+Ll7AtvMluxB2D/uvqVsB4e4D4ysWI
AMpmUziDtaLYLKC339jrCukbBO839HRtQqJUY31qKNaMwIxdcZZqaYjX+DfnGVqohS1KV7KmRie+
pgBl5ySFAe2Kce8QrFFiqdI0zPrzjO1bVfZxpTM8CcvjZR4fnfIaMCqSWLNVv5N24kNp1xZ//+Ej
snRyomxQkBdE+HPsWtX2IWHh2Q3hyVaNziaKVqpqzAOS6hBwrbMtpL2KZy8mxLZd3R+bl3lKy/NK
xBEDmJ2RWOqiPh4yJTRajMAmVLf82EYdEIFRIcKshFWA+c8KX6neLkQvqFSi1SNOkhCtofQTRmm8
NUYtVOSNQPCKAwb/YtZUykpilCs1svhoA0phOPqPHDqAW5yQQr5PJVoB9Ao+AHmlIWNzsQFjHZbz
ydpr599Xcd8xGkXPvgIKXN1uuGvJQNh/HZ0xlrgdfu2Y0QtkPhm09ixFZAs5WM7EkXXKnKOnuKuA
iEIjBvzEebSU+OrMT25rQQ+ifSoG0vizhl8N7DJciwkmx5VZQKkqhEyXMaTrCP+/tu71+57foaX6
qKpqZBH62346pGEnLiS0AAmqNqLacR0skFx75zTQHbshFlKuzqKhoT/G9SNtdPN/FjoyY90vYA98
WFmQ7lvUc9lpvlMTBkQal+ac0cFrhL/6jTnmINmPTslFafc05AWXlF/CgWxsLD8xtrpuyE1Xk0CT
ILpl1kiUoreENoLgd/eU+9UQwlF4P7dW6682rH3CZStFaeNOemyoKB8+KKZa0ikmTn2mxd76FxcU
vzPUjY3PfOz/Z+T4/KuS4WjqnSLATI8Fkcai7kwBoT812PyWnaMdxQHz9lJrfT0vK1i0Eo3Uiron
WP8/tN6zRhulClP4Orfw2Q19xWvLHBzwXsG3FJpMfiAsKTJqCrYTAwaWQSez7KnKZJdmt1LhBwhL
FyzAO5lGj0SHGAniWEgqvMU2HQ+kOTUuB9l5wq94x2FuAMxjLxNylFw+09UG4hsvrEdgaHIffL8g
t7oSINY2wStuSizahjVQayxWoXwkc8ZXSQci52BCV7sM5TnirpXKPjoKI/wMcaj+Ae+5ccDHq5CP
4LP8BOpCTd/JedxqhUYJcYmmqoQt2+4pCiu1ILkLWOuzP2hglnytci7cWKl1MiDGhRbYLu6Z4Ppm
+UHtguH9WDMBPFeWMFzP4aH/IxFtcvAiPDb9LnrT3sm3MZzuYaEmlQVSvADw/lDsspoMrW8PNIoX
okaIFgOszH+Hq+7+fhX/xqvQZvEF1PrIIFjy29JXbiB5U4zaa1fmUzgXk1AXvJwnwMqc3DgZe2EV
0PhuaTadwTiuzVMuDOcSmaquO1vGAXv1Kpn8LkK7qpX8YyaE3ACg8nqLw3jtxjirkXWrBHGXrEzU
g/5Ajyn/GDpVgPhOjKQpg8/3NJvqM+z3oAxVUx+jpFxTKymCkFdEerfU8FHqii6iZqqQ6sY1H5Ja
KkOjpN4veAJYa/ZPHjKzPqgmE4ESMGJxxBLBr79kdgiwZX9+x3a4DP5SazOcy8vz82w4q3imywjr
fUT2//yapa/ib+ZQ1h7sACARMUGDLVZ55+8+e8CBwZ6x6FHccZX/TtuEz5ITJ43T0Yge2w31771i
c8ZZRza5fRjzjGHGoWvJjQJeNI4Qx94rn0/fm/My2yqFp7sz/KpwchW8rlmSo8TQx7/AMjH1FM8D
0ldJLRkJxamentMwHpBq7JtzNaXgT29PGip9DecN+nF9HKbVz7DUB9lwpnOwCSZbbWvdrbkXouzv
M3EshMRMadciYk1vbvAuBifQrE5hbfjpD43Vp+V5b7TPXZdY4bQSK58JnIy5W+1qkI2TnHbNzQw6
Lheu/hFrTAWNGQ0+GyfK3VqKCH/rynQoC/hVjQmpsLpCkMQDSP3P6UDqDWzk+sQ24gQcshl0J631
D/lIONjSjt6Rk+RI7sYYmeKxyKtcpMnFN1YgfKgY1A25RzQGfwW5zN5P6sGztNnw2iTRb+L/2Az1
iRloCxLbDgpQhJw7GrJxNt+Oge7SHQbpx0Oh5GC1PTT2peC0rh28nDSyu6MJly5+Df6CrYt3W8E+
d7lvACGpPTN314BFbNZHCn+v4XsCCGfLjGqjMRYIE2HZgx9KQAX4fYFtfZIYQT0JI84BJlH2QZpk
6RffhfZdV/PYqZ0J8CT+Yw3B2bdrNlV2THRyvRLA0sq/zte+9SAsSpBQuqEByZKGvhc3Bo9qOY7x
bfd3VRhJgVGvkyaAFAOOs/vw4wS/DW7mmz/OpQEPw6mqDuoji4TQ3zu7zs3onS5WRZGgOZT957Pz
i0oMvzZnqmWiR29wat+7EoeBo0T+sBZMeK32gIJSgiGv1mgUmsSwVuKH6r0Qx2R7HYxuCChbe6nA
Y+JjuoBi7++kAZIO+UPjgx7+xZB1gp6mNFE9rEgs4zJzjsjeUlsM8ItoKbK6tOWKBjCd/dgGcm6O
zKmfhvjD2Xs2C0cpY4Cp0vZm1BXvUny/fM+jcSHGDx06aZlCC6oRoo/W/sgeW1aBfC20qjJ8DUno
GUYUrd2zCTnWrpsCgMhv8XETRaJ2Vy4xHpsP06Z9mfsP7R8MKLzqhYCxZ+pio02fNalVZ1YOVIzQ
iF3CbxCqle+ntM9MlcXqBBIQRweZs7v8ZJCl7rGXTFHMefqBJq3xOdbuvgovwB6c/noHYxqCaKRL
W49ihw0TSL3Ifo2/jcBJ+HPp1oci3qb71nUklXBJrRUHb4e8kR4rYyx50EVLQXi8myG6IjwIx63Q
BGnZxZ0SqvAtDx3zEK1LYjLu3q6PHqZwe8G/3hfLpUlXifbQRpnwwU5nVitZ2atrR2E65wl65cPL
Jk9vZiHjZIch2+YbTZ/io8NE6bm8W+xC8yoWF9VAOvpvzib6ABLq6ZcytXXnKfPVcoGnUJhbB9fL
7d6Ts9nFWYbBp2HXKhITPjsEwZaHzjjbXodUtLlvDKvTFxPcYq5iWSC7Q4I318pCj2ptLJJ/vUjn
sncw3wffPvYUusnfX/d6sQVl08kUiOCD73Nm5MzRmD3E7M8pzsnK5QDstV+pFkw5GoSFKkNfweaT
vqcYxZfGsHkET29J+z67qyLikmvoKF/WLWUGqeM8UR2tNrNQRJ5jI9PrkAA0P8e5xg0pe+SusDKX
fo4FJo6SkFwl+ZdvTRtEr2pVDruK5pidNUEbsKu1OSnXUh4HP0U3n9hfRs4SFcsLkxz0OBOr+1Ae
2q8Tu8Zairzrw7eSUQuYIOGI5sRanIxF5FVMD9NMNACPmeflENgs7s0APpwJCm9JYER/D2yCk5ug
VOKxTvnA/fbx8vwpJCv64LNdiFJqoQIv8+RNY9mQNWjEOSiR84pXLEUfoqFm1MkKWBoCOJYqlIYs
1hHNFoUc6Tr9J9D7TWTMi3In0PGuw8ouJv8gW73NmxWfTYDvHN7Ihree4FGpfuLpbioYDNBiLaUR
ycyCg+JzBViB+s3R2922fc+6tOlKGIjF2bhxpOFF5JD0CGHHKXuZA19/h0+lAQ6kFLUiLzhOuB4r
7aiOqTA1D4XnLUGoIYVURvQJoSXU8fAQtE1h0X/O9XZwTQBck452wdcSTAwIu8txbpiyRL/SkYHp
c+P1C3gUFR/7sOdryegIlo4erbC/ZyrZMTouLs9nr+1Us4f3HVM9Ps0zt0eWEt5IQ3Xh5CJaimGL
mt5SfTVdh7qHTqaDB0xptyHBF8nXPaXpz+wPWxsu+wjReySwHbrwVAF1EK8u4GUa23aCW7Dx8u07
grWh40cJuM2Bu3WqoT0jKOjHc9bPn6A3s7XFU23pykVGmnKFO52TzOIyTPfmP1yc8MgyjNEfkY1c
/0qjDn2zr/23L1MdwA6C4Rwfu3ABFVfBJA2eFqanu8hkrCcWrV0aPo5uputsfKoFqdQsAqo8elDx
roiUgiYziPKs6jclsu+WNslBgZ4amg6gUheL/gM5/IZJ2n1MCaEXZxeixSZxctwiATRMnH3+v+Uz
f4Hj6LITrKmffHy9xY+FIz3WQGLQy8zhFK2+7m+3gzM3CfBTSRDLKWk4ZVxQjv+p4H7eBx+pmgdP
UNAe4b2GEI78SQwsms6q1qZVO/e5Id/R/oVz1Z3Xu+dD3LQYTq1zllQdtLAhqW8Mp6db8Aix5ORu
Ka4bfWrVmkifGZO8hwvQnsI2gVZX1dL4DOgFmfzQZKSrWJLSFcRpM1tCiEichWIvWIf5oLHQSW9d
BFIx+/bZ4gXSjxywRT+Res2hjbhjlCSlEY9GiIXLHMCRlqGG3FyggbUeZxX/InLggQPnst9+h//D
9CZMYa6A1U97QTnpdoMxNInEF2EJA8dttaS/f61Itdve5cFW4xme++Sjpbgg2vzITfbG2YiZM+b+
Fdc2P2mHId2/1et7Pm/L5yiuoVRHdoz633ZzJgobl+7JjmV1trrAXQ/ToRsKyWE/kGHmzyd/HKXX
ahSsBFoocCr/th5SDUzR6bgJDvA6k90tJDO5qbKHZLWTqAcZJaDM/xWDTY70N9+rTwLHMSwdSgvN
6JYgdydh03axjkxeFrXqUKT4h7+b3NC9D67SuQmKd/+yRHxK45VhQ2u7aeVnTSW9FJplQGjf8BBy
zNJIfBJSTAfycpq1zU31oNu8vMc8cvZah9HeX91xw3L9T7EU8aU7ZrZ3pbgClOjPjC95Soih+9tV
UV8B3vpwFloowOuKkJ0Zvi5C6HzkgEltF3TC56AhlCVwDpsDwydMDVtC/g0QwV7biWSoxYF25Z7q
a7gxdk5m51KIILsCjxG5ddwm7Jk3jHiY7FsDhd6qmPcu5c+hLp/skxdRyAedc8qlRGLM3cljyi0+
48eIAUb3ubq09rvVr9UUdA3p2oGds7Bqhw9u0VOGocUXAOho50y4Ku30kno+0I7PRctguyziY4w1
3E0W7v4WewPlj3yhBKeG+fDVF267/+5frutg1VHcctztn6vgu3BhBMhAg5VD2KDCs8iFyldNt1WT
lxhuRJVtrgFPdOHV3lGpRLL8uGXVVYNhRNVrb316fDtIoZoTq6WodA3O76KVARCIj5i8EA5PBqVS
I+BNzbqQab+jDGA+A+W3oKiDsx1E2QLJK8JmX/hhuU5dikmXbSBn4fE0WELfzm1YLVAEnkfhuaJq
Kc7/F8iWZnLy8NK2zp8AZI/aqXEXMC/dW0RAXQvSj9pwZI9uS9sGbwvpZ2u0CVqH3KrlfVOJkle4
bF652WCrak4nIDhDuR7+k/lUcy2pLfPqfnWxGapqDr//2K+ssA0fR3XreNAGbJHTl8n2hwj1OzO1
qEkwiA8XKbeK2xCpZLjkOQ5V6SWa3NPgL8/gzPW8rOHaQhTFpuo3DtvhBBdYUaRQrFTL6ym+R+jB
Z5uGdC14RHWBQnl/p4c3VcdcEdmZKsIik/zOqgvI7t3tLUUcoCh4OwO4GVy3zAl3/I1iYlZmB+6x
Eh5n4OK4Ep1m7DwS0UlTRsJY07dnAOTIhSYVvM5RdmiPbOcOc+a79S1O2kvxnyxShV/reVS32oTT
bTMo5CgFEddh1/nz65YPKeBT8NtmtRGuiIPB7K9YAJaHKQLrXMWbBHTpNaWWphV99Ivv32749Rwe
gtiW7WLnA6NPokRiPRIjM9zEQVC15YLUrizAUXXC83gi7/0XJdNvxH/2Boa0SbH1wEFPk3nBTCLT
i75SdhdtJLAKMSuujVJEh1+/BRY0qGRL15yj1c6JsY/JKRH+6LMmlkcL73G1sQLNf3Z5WNrH5Zxk
KTIe1MnyuQkH4ggxSBlr+drq3mbbl11cbjLky6FrsDVwYfjhyILeFERAADI17u94ODn//Gqjfu7n
ItQDfgJBKQfMoKQ77MQvDDAb09qerxt7ajVjy/KLzmOE1LRiBhd2Zr1ytdjDQSV5d6DLuiTfpm+r
b7V4zfwOIuOGugiWB4DyQvblmwwe5KjS4yAu4Du92VUbde0catysDDRbv6hrQN4mIsMFCvgHhuNK
T54QzKXwaU3gFq4Jtzz3qkgLTGYS1/gskAlX7SzzcTQjYaa9jYi7inaBdi8rR5XW4ZjRQrVTfTso
Gs3AqluPGfhJ+FiJA0FdPVMZERPNELzPjhdzBVa0tTTZMqg+dUdbdp9B4gUz+NH4PD8sPO/q89Se
7w9DFgGr5/y2n0RpawKHF2UNQpYDWS5kp/nqVc3VrHiq/3qyN664yka45ANPrL/YRF32fOjEOWsv
a0RBx/gRsz3aiffQXgLXHK1nwf4NepxIF0gAgwO0yUbcnzDVMDTWWbPJ7/SOBmH1mizeMuKnV4jb
23wWOBJLKY4+329JYBb1JJwVwqQlwUs2o2MkGODudIIzGsX8WmKqZKtdMUm3JCbS4ww9HgrpC/V9
tIaUVwNaSQwkz7l6lkJUgz5d96bBY1N2VXn8oYf//VpGcGFQVJYg/rEypInIWqVtHo1nR3Z195nA
pQVJDUNtM/nHr/nZhPowWFOruRlo+A7ufA5VrfUKImU5blL5NCa7UuGpfru095doORyHmhs8RVip
2ygbFDG41/B76cODnnm7wR9Fq1S56kxCky89UoUCQ/ix/1NnnqWx3K38Dyj8XEePSWcAX7z9HUeF
YBq1wpzMkuKsWI92i+YgaeiCKbaWN/aFRkhMfbfbRBGOq95QpS9WxGJ0FpA53AmRxhWkHLXwqQtH
eD5IjoL0DGcspdiY46mi4fmm7DFayrxPMt7pniUqfU7vJQUb3pRhDto4b4ofdpgo2uCmfL3i6x05
obWyLM19CfHTBVBnjt3G8iX3NHCVlHgscQ2EM+j/jff36PPkgB1tEalmCjEor9PHFu02wwVoTkCZ
y4cg80VM7bwl3zpFpLk9S2MROW0quSA2n1G+maHb8icBi0zedtm/hGzEF5VfvePVX4IzqN8+DQjc
FcqT6S3Dyge4JCqmcAMTHJicUcyCAfx3IY/HLqbv56HzJCy4ofzVGahreByp92HrhuhWiYV/U/jp
ue+IYc9UjeggolyCCY8pFhji0e6Sv4CWQpHD+xLKuoIEcN4vnOVzRPRULVJy/0JINY9a1riw60tj
YE0tTKSy+WVMQ8gGovJqDYU2wydXppv854R5HcA+sNx/xHC9/vBrpUk2e8ZsfnZpNv41CYjTtcLJ
dGqtRxy5l/UNMlFyhZH9/wolLZ3T7XjKDNk503AaJLiAlh/ZoGeZLvVLRncWDyBNLyJ/JL0P2B8v
tGGDf9ABXpmDWZBTA/1DX6URLowDy9lUm4aQ3GODI/unVmkmjOxCE1iEMM9HEyQKhf3o50s/UQbr
2DMK00+scEubFXfXhCa+bnpK4V2wNCHZ5wAYxclqB9ojebVLcjELFqqCM398E14ChExdJAxzpvno
hjzGbdi78xwaE7u27BV1iNCF5xNVGRiWw6ZeO0jltBtgD81H6jLDrWivLTAi1sQozuAa3x4aTyWW
iL2RleYwuh+Nzp3m0R+8KRTLpdGY3Gx6/vOM8wyo8M0E75ho37t3xxIoc9vPvwDaU15aOW5fK1AZ
waMCBvl6emXbJoIKR+p+EMta1M2OpbomTHMWIe5FGxgV28UgUurLdLQki+FlvdjsEGDdeyTxTGoD
XoilrdgQd9TM0F5W03zCdmCOFht46k2peOL52kIZ/ypubBmkbhos8fgn3d6mydPAA+tYPl4mK2OI
RoQ5hStjhDmVkf60z80uIW0v4cP4sD7VZCKa7t/sCG7oIio5n/EzsnHztoJKmxCJooYgxGTIZLge
O4OiN7KFTRu0sYOhJD+wgJmHH54hiH8LRrS47w/On+2S4p9uxnlkVqq7zf88a4RU/Ff/1wScnlp4
EMSqwBmUDf2z3PYADa+Bn9YpTslAne39nr/OiJoWaV8mfqkhjZm4z/A7q83u90skUmj3vpY4clPZ
xagRegsQ2BI1N1QK28PMQxLAQ+q2nZDynDQZ1i3grXOuzraQ4T58/7Z1Z2t3JmmsJ90KBIWF2aTR
GmeapOMc7lUFaFCFKUxtOVcZG1Uw7HOJRcN6HJt6WdBFNq4kbD4b7Hx4WHashURU5uxLz9w/upSb
IycLxEcAomZ+O/cy8Kv23EsvNp0PccsYdzE3HCcA+y590I3TEgSv1RJPxiuu2CmwyT6Rsd+QCd4m
jtUwWb/+AK1tEO2zNtNPLFTrSTdvKIsteMmd2k8X75t+hroL+3LRwaSdxzYc+nklvLrrTwtTtozR
se72auJ58wUaqULMn6gijSuAbwhSaKX4cxjRmPVcDukVTLi2OHtHEdcojnfvPx7E0PQMKqChh0RF
uKcJsJ+T3CoIynN5akw5+1iJ6KzuTOQB8ebdl+jVBPunKxtu3DVVGC0cucJhBNtWpO3CO5JeCgiS
ZFMBu6uAT43WEjfK932TSlOQxf6G3iFjgvCw8b+7a1IIQjlX61yHD1DplFAxXQZ/DgIH+Ymk+yAS
EjAa620nnEnrDDv5eHs1Xrt7UIczx/IVK9IhTU0kWgwh6MMRhQjnRolh+WKnCwdih5zJbFcZnVpu
8E7cwL7jrqrkt01ADjHomCud4thNUWxwcKEZMt07BovJTruXt1LGum5EOfirOo/VKzwmzkKMSDcG
PrWjVyLd1mQgvRRalDMq5cOmWj3pCVRWFrVhUCy5PfzZUAWDoU2ovQ2bjGevWUV2M42qKkTFrwvT
UTu92i5eynJuKd/VJN6ZhvUQs+KCJJ9Joo3Mqblhpxiblt0pDRg0MYS26e56++P+5AEE3PbRVMJp
TPUJ/JRNEyjJcfDZdUT82Yv2Ydc1lQSrMpELCelNmyGuGggEWaOBly98oI9fjmEwaRPWlbN8U0T/
vnX2Geay5XgeDJzE9joOmxR85DM3odJEHfiGDCqLiSvmeivHwheLC7TFOkIlepRrqxi3QUGdIuIq
/kDej5YmWtw92l7P/ZRLGrGEw1LdOTpPTVDFvzYF3ogxnWNr+F1fixRJfL3DF1Bq/HWD8pdhQtkZ
Fl1BCUIoNc51aECAiexgmqmhFqZWkgEzpkQ1mq920gnzyT1FQlV6X1GY9hLkWIUwkGlRjfrsLGn5
+rYZSJNg6aAZPQPoBGMra1VeIF8bl4b1b0QEc9TIBtHGLJ2HBlpXwAkUVLyHx/tTBGOLE84YIOzN
kltQX1RmwwySpeAtXKCS09KgkzWdRQvdndxD2VhPqS5N6xGJ4xlN72CGt/9h9sYYeZxp8bVqYvdU
9JxLY76VlfOQvroVbGGvONYkN99uCC3ZN4/LOyIxlpDRW2UV8QvMGYJPIkCVzlv+Du/VYQt1tbCM
0jde+/nuzrefZUCGqyfBR/iKts/f19sxeEa4gP/qmNZ7dcIYTUbLcxfmRu6YwTgPpE2KE0vpJTkY
F2+PB7Xb94eeIH09PB0tuEA9CygI/Kaf1Tiozl02j6Eh3VDWtnwyYFLYKeL2vmI5QG8xrBL8RhaF
7UXNUcOp59BP4Lx/91SvouEjrBcp+VhPrwgnhbGkVnpEzEqMNSRP9UQGz+NWU9TZvsdfpRhQ5g9C
OyUdLDdU0SVuporoqNWC0mvzl1CJU37v0F1YHQvrzokjdGfSaAbtcJCUgGKwoenRwyjvVTQuLCyY
IkW10OaJxE0Q9PhUDVZwTsyzYhNIWkZTBae1oZsvXlyuVXwJA1QeU3NEA8P/lK/75p4o9rCJIpN8
J5vl3FFM9L18nv6HNmtyhl66Sky9btaN4ZqL3IvliE9buMegin8jPm4KKVag5P5/qNR+0vI03kd8
2/p8jrjnDwsSjwju4kkDpquhutFGEmfIf7Qmv9VLV7LsYX4sNgjYFA/+VPMgNy6fbSgGJrj4y6vp
4PWMJJZTKpBunLnBgCluFv7O/FLF6AilPhUTNyzvlki7QGkOnoabrfkYf7lCirhJYp0R1WyMzi8z
ds7yqvv/gLIg68eVd/3akqEhMgFrRiTTEvXWw/JJyQ1ff/eFt+HU4WfaLn+C9LNJIYt+tCjppuk5
7Rfiw0dbYNpwPDHo2DLTATiteppsXLt5wSYTiv8tgtKyempdiTUjcE+vHjvAENyLiKfMArVUzWtr
5pULfliEiPgkgYUFK8587PB7/6jamG2Quu7Yg5plW2lr67CyE+soNSrwCrZg8FLW0JQUUALUzdxh
+fR2g7/EPwmJV7+G1RCbr5223GGTY9ntuiYxj6QNw61xUloGq0qIZDkkMHcMlX/37jbeZkTSrIpA
6K0+/ggggY7Gu5V1D2Py2PapSvcxQYkGAbptGakJNjjxiPOcQfhewQm0gZPSBaup8ByLJIzciT4k
4z9H7J4aOVFofbFG+k+jCpNAn3TkZfzY3+QHKkk6E5QKZtN35E7NidXePuIuUegweoFhPRbx3mbK
BBvG/70cU/g2QySWI6eD/DuFDVKXlEY/wxXG5d5/udc9DarCwMYa080b9TX2I3WGlNNBEyw4nZFX
CBoop/Q5z+IDTDXOSsquRLDtzWHkN7pguFTcphLJm5LnWZjyBSDNfN6wOcn0ppImExnziM8xJpn3
ayJ1Nx4j9AvByz22hHxcgzYLmoOys/kM7sF5dXxB6fKm/EfWrEFhFH5tlIY+ElaE34OSG//CMEN/
lSLPpJduOsLLK72R+UKJ2/6GohR4JZgXhYsvEtVBtaiiaR9lPB4vg6dNfYlJuLVVq1cNQf40EPZO
HgRIMYlPnmNMc41F2ORKUipfAm2+MO3IvZu7k47cNWPHBAHN73Cv2TKzfYjymqsTTtI6VdFN6x7R
qxnebEQ9ecddbCvp6CxEdYW0Dt46pvXVVSFsRsHjuDMl5oFk4a6P+tWAxLhrWKoSwYjdEV5TVZ2B
s08Uk4TgznDDqN2RtNmgJJ3lmkpfXms9tojC/SRbg5x5bmSGdEupVEh3mMuIEGUdAYj8RpBdLhHx
Hy5TXtMgWkNK/CzQMBdSugxTfBoHSubrb6U0OcI7LcXqSCYIXYuwAstoQwcojfM1y7VrFrXjW3Dn
rxQT9jSvM4GLQf87A8VEA0toHDKm0A5j2xvPHEyi9u5n8uW8d4vLBT1RfkyQm1RXIvZ8vyV05idF
tSJw5H1WOfMbu0PTaXMf8jaGNZxFhapiEy+Z466NvLnhMwxxQ5EtKulQjI44Lj9DiqVWklhTJGAh
6wqzM5yrjRuovvcRheTq5LStBlOc0hQffioqWgSdKqgBZS9JhNdgk85rnugEAGCYXgovoVPRtZIo
Kt34EpNrffxPyoh92GVUZNpm/gCb9kS7QFSZj2UDMArFZpj+OdaAZB+Ol7Tk8DPOPbXpzsKRGbWF
i5YGTI7jHyYu13oKdffX3VvxClCi3xNcjobuvWCl4QBYFt+g0iOK/jNWSPlulib0WraE4rogvLii
xpznmzEFD+7jXe+hMO2TVcrt4FFMZZvo8MQSCqh+vKvEeFjSc1ZVTU/wHYQlbY540GovVOx4Y1gV
h5jfV34lsmAOo20VDF7Qzk250qTKbFsh4In8XzdatvTq3j29OCXtgXOVGvJIV/s9mvPhc0I8WnHg
j/ih85g1jet2KyDZY9RMq1w9PFbIUSLnJHT4d0ih4k7Cr8jXf6O/6Y/MckH6UBKgkUWAX5YG1cfn
pb8to03tyrBMYY+oCvsYZnZkSB9U30ihTjGHlFdxV7E5gf4yyBzCk/PsBD3mz9uhe3ap3hb3xuVR
uoFgESf2/i5uTFAaoqMqwfuH9+thLZmM3Z+5d6VTCduVeJSwHlH7V8m7LS4xAA0LF+7sM1R2hTY7
BcLuzRcSgnNfZHZRZXYweQi1u9AqRuOhVXAsEBjiQRX/iJ+B+9HeYRqYNgtRA/WW6o1KDZv1fJuZ
iJrQYatL57B6JVZj14A4/3TjN1b1pjXShiCrG1m1O53wfvzpDQwf3QKlKTa+aOimTFC+aIhcBZuj
IP3xfpsF4rT22/Q172cdAFVPLOZX1UBOZOcUKiBWYMCQtbmfBdxgP2RwBSU3rrKRPQr3W2xXIfQ+
GtXOpBjM+QLVipIbFIovKQpRWH7cez60ZlAnzXiwvqlfHw5D+6gPWsBJxxxKuECDFwAfk3uD577E
VbGoQPBxUbJelCtXm0+dJeZFhdjckJ9iaYc/9Ge1yC+TQREK+OQdl6j+ZEBoTWVN4/k1PB8hgPut
IKXKyhJq4FBd8nPNnTYB6FWo3SExvt3Ya/I6Zvf8BEN2z5XcJJnE3j56cRsjP9YK64zMt/+qkwRk
PZm5v4L4OJvdzBNlUQXuk+yNAgCyYZvXp1XvFH8XMnTlFZMYp/w/1aDhNDidE4cqwFGprT3fhrXi
gnYYiSHLNmdlsHv6a1COgP5UbRYaYmwdW5GHIH7qgbSVgHmWkRnQDj8JEnkk8YcbXZZ7zQmNssZW
bI6TJwcpP07Bgr+/Q3fR401yOW1ejDbVFjBRRSwfltjMsWp48aAChVBWhUkwxcIhPMA7NTZX+rbH
sWyK6QJIfgqYZ18RdvfUjQBCedSoGuE6CSg7yqsV4O6vJ6FVqgSSzFY7H9gdsbENw49MmacOlUjq
JclFV0AHRm/WPHOhjI9A8WCq+I9G8jSrZchpDXqcyqp76W/1YkPBeDAWrzghJTAJBsnVc28WP+be
HTPXoSoFcYOfmo519eZ8s3qxzKkPVjX2U95nBEL4TEtvcL56Fm4KgbnllN3C20ug+8VdgQ2yr1D4
cLp87ylhGUwR8PxlfWsHPLc1SM3jg/SVa0ZORpPcCdAWeHcNwRoJDFqZe0/lC/OSPe4CFz4420pf
uT1mlJV+/+a7vPD0WMeeXGI3CA/xvgxmaMJBvvg02SsfiVz5hwTUSVefDnJOERTm9XTZPcA+d8m/
CoSD3Jy/dHvQaIwa4869Z6KTrQJxCcRcjl9eappPynhFvJgHF+FvyAQBvoSXK/BcV/+oZMl2jwiQ
hae6iOECp6WA4wXXJKSX7ko8eUNwe0yfXW12IqdMnDQ3DZ3z4xbQdMfcGmMvHKsZMEWJQq8/wDX/
q+4MB9+n3PyWu1LFDx6QPkoNT8LKj4rcN97vzbMRHcfO4L+GEQypOumLTaCDPHx+tTmnh5kTu4Lf
rULe33vG/QPGoz/W0uwEBw2aclY8N04HVKhrrkincx3KlHDUnEK+sL7CoLDKwGUHbE4HhNgbI+HZ
U/qXaQ7JG+KT1FNDHkw7PNkZlzAXwqvablNfD8HORHdKz3DaInobg3gutWHRevZ9ixE8u9whqa+i
f52vkrQcMoVVTqW/xhHN98zTIGgTVORHbTspCmuQz/WMpO3yHPRCZ0vGsc/NUVU5+HXdrCGq9Vbo
mmC6Kf8+DzpY5ynLYR1v0lQ26nL4+1Su+GMTbhsMOERg+Zr+T8xK0j/yRHic/ITvAOZv91/iXvOm
nm/Dq7reOIeTjXIiM74YnIpmLv4odgHp7Ff7hPmmD2e+YltRyqnjBNRuH1c2jh3urhwrdeG4O0SR
3QAVuwe4TINr18AQrOSlaYH+cbMkk7KvWeomnVJQ7XNY7Kmx22psqIzXjNFIwDukBXuVgnFBINhJ
tBZGT/MsoZVUh4W0DWorPqMpqUPyab5n2svuutNzCg/dP/OMUO8nTCCS2hkipL5yxJdxYMnWhEvD
sVhg5Sxt/YpGwSvtH11jcEgb1/BpKmyBTXpcRmuXtw8saUQLWQSeTUpL17TLPELnS9rHWqbQ/MJs
lIjAtTFiEBe1AgEuadCiMlRxDIPmbtjZ1TELIlTR8zvGSPKQcgGk7E4BXYBGINJp0jqKMPjtlpDA
0OoOLZg8kHQ5oU/qHwMjrOFsAjJ41UoG5aVzuaSkIu/lGISmmPuFlwKor/Y3Z//15rqBJGuRLQgS
DYTx1qcsgkoHwMwvadXnGCz2OTX5KDA09oSocyQ5sRn1rxqd1zdd8bhn2OJDm4PkOCDJqotTEdvt
tXh15xaUTKvj8VLlJkVTan5B6TmvKHAZbEYx7XR7idg/FJTsl48daTzrOYC1V6TjfqYnvNSRpqvZ
BcmMlawwT0rrXKeRVvX7nteZRE9reqXwTBEcuTTF9DWmX0pHtr7mc4ERR1Vmd7qglifRKn+hNVio
bSvdIvkne7+hTEoDYElLpl2fkHj0tXrp7t4M5GlqGFPj2B45g7LEZWi6ymYad9fZd/z0s4ItwcjG
Cp+EJaT13ZxyEQJm7zKAYi2AOSqfDsnZ+1pJH0TobkDmoFc1Wok5C69s+BA3VcRPJz7jWLWwz9gu
kypZByaltMYAqTEQEci0OHEPZWyzwGO22U8DbxFpqQJtgkRwtGXS4+hVDC1BnJMaIYiLtDWwBT/9
Gifl508coeIggJYRQEU2YJ8hUEwuOehEI6yhf401colZKjQmmRVpuWsV5IA0Fv9ZkzpQAzPSy4Z3
3xIRme40ylFO02V+AJN5OmI39Lv/MM67NXdBHcbUC2EB8rzzTA0MgL+48p4VCNo+6Ihp6eITgvw8
EOSGzTnYm6Q+nilnr8d9eXbFYfqFrPjSx/fKrVH9GEcTlzr+GRdKOdAdTy/f7LStkaHjOOvK7XOg
xSJdqyn6v/IUV/2ypHNO/r4qMvMDcRZcbJ21Xc7KJgXMlzket0hXKn0eqmb30myL43uFQUgxdiR6
h2afHduDaAmvC4dgD28he5wlkAYl/paVsX2Gm9jfMd7O9yE68UmwWv8IpFqdJqpBOhf2q/ObQxJr
G023D1qxQ0SJgAsZirKLlyiEYYEONeU+jBYUzEkDFjkg8Xqd++fQwb8cHH67CkVWIf3Oh8GkwqCQ
EhTIxZgdyW1LiQW0M4hjKF6pI++LBmPsE3ipWhnm86K1TNsJ9N8++08CNHPh8Uuv/XKQCksnKPQ8
2cZAkKCALkEWp9URr8pOzrLXeRcuAr8ymIbwMCq57ZPGot8XzQKP2Bld3Li3WIPDrnREl5XV1dPM
tyoKgHSFgVT5XtXUjV6gk1sqMnYXdcU5d9DA78rdhfH5iE8L4ltytXTI0jAPQTQ2X+Pyj7JqgukY
1DQaNynPhMVcTmdDfc/P1F6C5CNlSwn78WDfdtwKu+GxlDe+YOiGVKPZtjMS3ln517yCLZ9C/NYx
3I9pO3O4MPgwTDK/AABoIrTz3+DZqwxEljUcYmzi05UJxIB1YsY9PZ1RhEWp8EZ0x22HfaI3IaSA
Vgfyx1d0bkrIcrMZVi9fWferWEITzsm72yFGwaoLEu58wymDBAJj8i9AZBt+0WBcR1X5iX07jXkb
t4brq8R0DJCbPfZDJN6a9I65nhPZcTlH6YJ2hOf4V1+BKzwujMl+44m4cyqtyrLTfnd/5g+7SY7i
c/WxGcRB7aoJAn6jXSpVklmyGrPa5EBXlIyEaimfcJDFZ813vTBVVXmBpwKGqsSZ2Ykls+BZOgqz
tu0lnKYm7WWnFvM8fJl46WNrU40cSRa1wGav2No6z14c3cmBUSqHg5luxgPfwa/Gr5BWE491+5VB
difX9lkqgaqOpqk9mGw1NcqHHUFtWshhfj6Bt5V0IMNsogTsdRmF1UgAF9lY3XUFf7jByHCv7bjA
BcxM4+GWy+zcuDWX0lRofJichfCgLrtaHFRB5O4g0w2u+kHdcV9GsEYavrDl1tUht7X8ugIsq/7w
7789nFa0W502QQwf6bdyF5rlJe68FFNjJZGjAMx5Yh3d/pam2Gl+Ukd/6NdCymHaHr4Uh/lpYmEs
McSn5wrz9L26OTSl/o4+d5BgSVmfSfMK8s3d9Bxtimrmw97/+HNh1Gmpc+4vSjbAIRb1ux+evvFO
KFYqD31P8XyHyvfHMTo3ZLM3o2q03/n521duBrQn7KwO8mxN1CkY0rIZF22wRvDQmmdL6COW7i6n
Gl8xEeyQU4SA5y1jnc7EqmiHKectH+6z70Ule1mY3nFS0BkPSrXD8AQ1nfHZs2IlFpAiYkD+3rKe
PKXiTKRhn2ivN0hEk+ojNhQFCvivyEiS7vJLYMEwDiZZYfz+fNVXNPku41Pc4PYnohl3DWIyouTE
pNzgAg/vzcXhNc2oMU9QprkWds6ALwVAGE7mpNENBJEdgMN/Yn40P+iG4UsI43fBvUNlWV9oOQpq
dXIqMjuT5ZWUrqHfMgJp/LWbEjwGvVKDMvIQkrKkazmE4Z/PMzOLd7s4DqWKjj37ZFHzlZrJSc7c
EhWQSNeKRcZ92ANYUYl6fF68p0lttBXYhGD2MJmjRwbz2UgTzS7pfIuN/XSleal9gguuL9zT+8tO
9oVYHkl8Hh8cxYGuMA0o4BV6mczf/8kdMzOgt21agAMTwXggpMXX7SmdxcmjL50E0ZRSq/99qH28
cD7k4XGNdRIXpwQtfA925Lc1CAH7aW46wRv1AOB7dcP5t/rZyC15w3jMyWm+fAAhvkRPBShqnDEz
TCcHOrJS5xiy6IAUJB7m++CU+0LgPALQ+/GCgjg9ecRqkYtb1EYUPIMfDKjsGWYvlXkBtWKMuUyU
lBPCKdL8sSpJghZbrtJDGHzWBPKg/dIxMFjXQctGxxbGYOPVrTyLw1ssR0IGWQo/L9blC3pJQSsl
ZAyiFCFfdylFhP/aJ3jp184/Ic2zb5QVr2R9y0jcJYjXOH7FbLKlKqYvpkenSDyoJIl7kUXWtLjB
AdgcOuQAW7ffFNBQHwsSbpfTmyOl7qVYfkayHqSMl5zQ3lGp9hM0yTgk+BK92woRMUe833jRsY3m
dh9V7CkQoZSqzw8beBuMndZ2UdrnJF6P/dGKsrV8tMOm7aV7HNA4ecz/kZuVgwHAg1OwbH11bprf
Qg7fLzgYlCxRITYpyMuVp0j85SDlJiwojqV9oB1NTBU6L8M5O9Tfdm5YUfS++g0vCs7cIn3l7tMi
Bc0cNKHIRQM+/fsbLQeF0J6oKdx0ZVkr1aWwfTuM5w+NDolxjVW4O8zbqQP077FuKV3yS3bLPp9j
HxGtLh+mvZ2r943c0LJYtyfAi8awIJ39cW49s/WNyn9F5Cb0W0YMgqguHSkxSeVHzC51YrGiyPDX
8N4te2gADbJNl6xGbfeVRW7gb85Z+fDoM1RTw6jyeXKQNCu0nhnxet62f424hO1uo/i2sM6c8gpW
oMLluWLaPqj01/ObSLar1j3KsUCfYbEidzNHhIu3IrZbMkSw/7mVIdjk6Uano+qi2lh6epHjDN5k
9VOsXyr6MzZBl0/yPIAZvViFUBDFOWtYvi8jSw4zzaYHWgVF8Du+XuKVzJktEKIL/a413nTILsEt
5jtdd8Nr49hMI3trI0u1dXcUelsqO5F7v5jdGnvpLKDRMplnCPsDavuXEtTAZXST+6sToVllnk7z
yyWl4roTP6HsrjOAX0RC24vU7GCPDjucnqrGd51+W+i1jKUqSftZ+dkDN+z7TqzX0j+J1xjTk0s5
Av3+KJUyRqPx2flVVJSkPO0Xn9lE3FyfXTEe4+FNMKb6TAKRNcBIGRi00ZKM2X2TQFfB5utv9wnI
fBgh0cApohX/05SqPEg1fF1ur7UBYwv34LgK/4nw8rs+ULxK846qJMBwyQA0BxDVQJWwkTIw0P5T
yU95PtB4K1fkG9Sxw49H3eXMJb4k16qjeCGDnpSxgFeF7/FyDl1sozdiGc/d47jKrI6/8zPoLwpn
cYTd7o4NQSraMyqNdGkn7ayCMzBeJ+cD5NQdJIBW1fBGsyScLZ4P/MKqNHeAQze5N7PSxws+t4t7
t/x+HztUaO+Zg8FvjRej5tYx6qBFQc0cozD3gqg+larv2iuIR2+eKbqnl80ZvuIC0SM/cWNS2Sb5
9TXEZNj0iaGGamnehzM6A4+o3jH9di1RNhahzBT2si6WiMC8+3QQn+dEgWEOG2xYdc98ZNjMsqeg
fMPCSIDTRVEVoS72+Xt4Je8S9zWVpfXNKrMN7TVXyM4n8Jbvjb9x+BE+2exBIt2PM+2y4lPkang2
waYKk5PeW8VmxS/zLmoS7qIxgRgnddQfoNp0zAtFQQxpvHvWrIEoCioqFJIYR7SGF2UIAdNVw3Tv
jOh1W3Wil5OEh2GhMYi8NAz8zQOtYI7jyrJ9wDuu7a96qkOrQPAkhNaT+1qA56JIu1wLtj4U+4pZ
fX+paw3uZtOIKBunE192PgUt9mQRc1UV4YJRHPVHasvt4QH+/xTIYuNf09omw++htsb7qj7r0FyT
HdDiIeSZCy21fy7/UYSBwyQs4ZxDCmSF4WJflgT2gkU2+Lxvdfi1FHGwjWXP1wJDlqykNznRb74I
r/KqNLU0rS5CIZnT89StWaq9DkQqfNsEwrHCq5xsfFtrpFUNHCBoH1OYf1C8psJM11m77JBVrX1q
Le4JdD5m+95tQc9+4itEDAowD0crvu77VdfgWgGiz9PdX/qmVgUEAHplSU9jDLtHSFOzm6QGB1jE
14xrJ+nzkAysPTDEk8OegMtX2FUg7U/eV6ClrBrdSy6QOrh4J3EYjYz9npUPUEgqnZVzBgIXvWsh
pTJpUE6frRD/96fyYnSbWhpR/sSOY1+gP+DpVhp12shGLlC7wBh2dNNYDw4/kPzdAJPBikV/8QiG
oHWO51f06XypENMJAI6O3MfKwywLKfkDkJ8iYQhDX6UX44agLGs9ir/xk30gLzNPeX9KA9g7zv63
azlm99uu2573zIFLECS6x0sbtEI+5wMDMkAbSjLm1etYaXcJ6ONrgYwNEIsn/QvJIS4L3x/U2DL6
LyYW+G8Uo7Tv/6vxLKg68cIfNtjadPDvLqSW5/X3E1VhSt6MIrzyAfLsTtLkhQwty11p1DHXsnf3
0vPP2UyrI7K/9Quz+rQWm1Oayc49kO2bC+k4cL7E0gvCsy/mfauruE8t9rD7+Y9asXSKigyuhNQp
D6zawpKSnS7ytHzenqvb7/pKpaT/d9+eKZ3p0YaA23yk49sHMbPfSv101q0uTF+K48YIkaFp9c6G
CZutKEtTSGwuMiPzxla0fTYktVDS9OJevosoCrnEe9v2Q/4Qo+v7hfL8bUg4UMeQW5f/vh/NkEgy
TCHtadnpzyUjHMQmmnB/9GBlZFfj839nulWQDwM1C5kUjTwuRCSeOY5ac1zX0ER3dIUsx8W6cmCh
cGzPXWDS3J2mVHg2ELTNP45L0GyDI/vYHWA+3rDu2ZoHIzerXqnX4bL6uay5O0xGQq27IKCYmJm+
NKzZ1AqQSpLnJT/ypHXvcWcfbOWstCygz11qjNJMhmNEyTYD8rfahD33qI9AKf7j5M3mIQ+I9Aqi
p7h3eOzRN2C8BwT3SConZeZrP3R1EyEkPtkFbmSdWZFGYDbH1O0meXE/pwnXbbxAn9dbRQj/9EWW
81I3YhBy/HKRDMYQqDwuPwffLEILn/AHuDOiRlPqEv9IdZOjxLLkPpj7yTRRlUKByPPQ7Wd1mysr
vULcQDjJW3U1sc8QRDV28vkca7e01L/D5AKZv/qTVRi5marwcu2Uo+i7qZ/XBQ2VfmZxst2NoOs5
UCD3XoUbd5lAtjAICWrFLKl9R2ixuR35rkLQdJ5hqDU56g7KPB+nqermoMIKBU0XCUXSeM1vmIlM
G0eZmAiaqq4zEJfEf1DQkLOfF1eelOS1/E4+lfKXw9WOYWeQROwUozTKJ4YKsilv2VqZyGb0nW9J
GTSzsSATZF/CPgbphLE+Om3jlvqG8ejfwxaycWBvqtYqYUPJir3kKW7A+FKfgBM0W6yQMdVYzKMh
tCg0MaOkRd9QgCMqz+PfJytLRzq9s5ULnl5itJQ/m50vwpU76s+i8B1CEByqH1Agw2z66YNxYdlK
Mrb9PIqq2C3CVG5aL13n8B/DUYgtqeP8VSlUyZ9wESpsB7f7khnfHLCbol9yBzx3k27VQzjhQTdT
ir3sRS3KM9uN7cQHhPm3Zf8Y5O9Y85jLUjfxe2d3Y30SbXSvAtgEsG7GPlVbFgk8H0FS//1BNAI5
0YmGrsXjIexTcqqtIKTxQfmMPB0vXQY3Rky3gQ5mj25OoUYhARs/X8pi/kcLCqMYAbbqDbxhWL6J
GMDSM9EHlYE+CNILqBMk7bNfP3kUO/U3FYfnbqOf5B9Y8wKi9RNRBuPsvCtj6BJkCu9SSpeQ6GEF
OIB84h/buB48WfFtV+rC9gnplRFdAC/pMNca9plkD1Tiav+I8yzDrrbdvEHBly1EJbtS97X5z7qJ
Qfv3DrFvrjIvH+yah7zdWl1qDZkBkJBYpHFQN3xlMoEToCpwuB3j8FxchIp/+W0tIH3YKl3UwgQY
NK+I+6jnmZe0R2ych7d6OXPOYjfDvHtdWVvXX/SoToY2L7O1PRMVnr/dLP/if7DeyLbkZ627ngBB
FcUq35s41Hi3ThcWDFTHHu8OACr5yTuwU74jahlcsszhbtbMlcumvtWXm37hieh1i8d+FzR+i1Q1
CMfFyJHzSoH9qCbLdDGzWzZm0s/lCZyCuqurEZQuQ7crdB3FXn53A96RPVywZLM8bu7VB1fL1kGJ
ZrMr+JVapLWXaygz5289+05DbC77YeyMEOlmKEGAIkjTC1kaWpauaESkxqCrS4WhPBtxipaBF+z1
4L1NcHGJ/U8h1uzOx0HBV6z2nkGYm3n3waoqi4+X/6CjiTaxw+6lr7OsTSM3e0E1KRCv5QtpniUu
M8OuzFKnojvST/3QnhYW4EqHGEGL/kpxGIla4D1LtMt48/s+pIqEa1dRpWSu6ONuSbwBvvrtCvyw
Thspoph70P/YaJf6XeqzqbORuq/zeJido7q97ym4qCavD0wgz72209wezOzz8m2+D56NvcLdUCJV
drhrQlrU1PTQi896LJNbtUrr64wcRFTro73gtmzHhWvxdetcWC3dytNiduvnuZT6605Yh9Uy2CEd
kTKzBahstIFcLLFoanfIS5wv54el+/hbymS7wdwmFKymk9+Ukym6IgTdsXBbBRPARZNZaI8wwhSd
PzR5XnUzEXGTNekgKyvQ6BK9EkgpsxoWAAsqzmaWKLDDgpOzVFmsPzSP5Wmbt1lZPrpnVwuSigtx
AK2RZs41dOFdrCxw6l2tlUx9+m9/U545DGD2BeGwHTBxYoQFG3+Z3sU0oAk9q4XeLRqlflAHajPI
4/W1M1GNLVjU53DN5h5Ors+L0WqJIW3CuaMIvsYbkW/JDpGtLAyFDIXMCnHL91SXJBib1n/LayK3
TzKiyfC3tRebGaMTbrsD91bUmu71vt7S0wRw3rJROY1Zi3z49UIBg6WzQaXbsnGE2TCd9gcgul+9
8tbkxOv4CCfIsMTNgVjdtyX9uwc3oewWgQJ3s3jTcuaITFutbREqk8kdATnnoPgJXWgpgU5x2P/h
ecp2CgSsc+OwKWl8PndlVuHj/vBgF0lDcJ1/TIMM7WU5YHZ6te0OXP8tmp9WYjPuNn6yOoOfbZll
DYdY77+AAaFmJNbsM5m0OAuMSH7LQMJOM3GKx4JAOtTWCi6RrUJjthScEjeneIoPYqqx6kVBoMJx
GTk79Oojysox8iYntuAl+udW7/XYXq/yStG7F3GOp1o/PHrKTgOEJLi9iEtm4yiHqCwYRh3Dkjzb
b8lacE2caAtfBoqtowkLAaup/GdfDUBlCkgs/097H4qze13boOM+onVb4ZVHJ/Ka2cd7e+QvJWPV
NWZkpa/eTzptC1b+03kJRGsqgT1rooGFAn2Tq9cEJjx3b7xeUihBI4LZ8ouRmaEjk6N38V4dpQT8
DujYL+PNjB2hXcK3POPxW6Xl8G4aNtNLjiL4+y2+++YTadMs4B8xi41Uo6ftz1W+NeDmA6DbkKtz
BcltgzHin8VSdcXxIj3qkWRIxMTC1MnOm0c4QUqpuvFc/yuuhFF9t3t9hP9aQWKVh2aIXB4tHw06
Qpm+Va00mYdomX8C0TPT27Io1AOb8ikLoragfalQUcfEuD1ejtdlgkkfkwdTh7cnaORuU0d7SqkT
Gc60dtVOgkXuNcESb8TJh1uWVepkgbbY3cqZH2nd/QvxHTNc7n4ZllHzSlpQNmxBoDC/PCjEYLbZ
8Jv67lPZCRP2K8x+EhSJePf8sOpQUKr1JBVAjHF5h5e3/cHZFKTzKp3NfiZ2Y7hE6W+sloDgO50m
H1+XH4xCT8w3gVOJWICupZ53yOCUl6+ykKsR3ktTEGIwydB9T6irt/dtCd+N/WgBKHKUUMWYbTNx
nEKDr+Tq8EIhQhflSxG2ggeuhr3o98UsrWsrYDpVuNmP4QO7yYwIyJVvdXlrsA39D2gB1KfNXrQf
4eNea1WLlNVRwmKTjb16B40Qn1RJAfrUAGe87yE0Dp4LWXtjGgGpryM7SuVRHO9rUebdLtDFVdnO
5DcgXL6t3JSu1AVdfMCgoBYVF+KInFtnmU5OKusdSnn0CSyEn9WHdiQlNgB9/PsLezm9ODE+m5Jk
xRKx07yTO4cK4A/2ZKL8Rh5gxv1B24OzMnJ2bxcI1YsnNOx8Sjga/ZtPnbj0+A3piVZ0S2Kab9iz
tyaGxRLnpmj1uKojZ/MIJHzLpuKMwXH8jMsYmxWv5qxlDdg+dMR2kAAVSRO6xe4H3MJbh+K+eDFG
2/ssDJeOeiLrrzM537D29UcUYtmZlCLPWudPPJZ87L5aEi0qxJDZu4IeicL7sOY9Rjrs7arYRGGp
pSm2P3dn79SQs1cBnMt/njWbKfPcXuTRxZq3cyBd64RZ2SK3+Q9Av1n+OvHBDzvyM9QqCnl6eyA8
N+GSC2/ZvmV4eM1bztcNqFco4QC1Sv4ILeWgoiIo8YsDsqqupjhJjIqzcFB35nT0EKGAFKCwYstG
eojfqi9d+NZzxx05dimap4AjKFOGztqRinMZVXhE0nHLn51T09K3z82ji96o/n3WurEPqS3oE7wU
NTwFiBudHKXWWq4KQFTp5tGk6SBcKcjnpYBwAEyCpo4IHuouRClxJ2/OJym44hP1l1K8Gqeat1Vr
UjuBR0/RAe26uLRr9g0y6o1SkHJ5GfOrHlmO8HXkvX7DgOQoVAvrkRKH6Qmiv6llM5ouHWijEg1d
56SFErwVg3ps0xr1bMET7TYx4t+31OcejUNOxxvFDj8hO3V+jCgfiPPzzkLve9LWXGYB4gDXzNPX
OSZRYSshjwqGLmvCo+qHyh8IpT/9AJ/Iz9m8KvIzXwCRL9pJBAkypEtbAMLHWditLOye+IGJwRsC
ZUafgOzOjqEHHEqIV00ezwmY339XPxP3Br38WFmVNfb8KkEgubDPnGKFiS2ltZ8o7HAFWtkCIIMW
s+huI+K4FZ6wMt4fAc5aYZLB3dWYcxOjxO51WGPkhbtzfTdsET5HOpYg9WUmMXO7rXtG7k/xIrBG
o50OW2hhqQYBvoCVEEjSRSuvqL6CXhJpyRclwBXNiKnva/lyl28KhHdcn/1fh76+Oh+0oCMHT+ao
Z/0rDmMrpppOhKxoV6smbOyxgD082LcawsKC6Ma7qrTSXNs4KD1yBfutzZB5Vrz89IIlbmFR7q1Y
uiqwBruzCrJ15O0xqYGeRIicmcOt6fKNXHBKkQ2BoM0gicAFywuG/MV7A50K6PM/2yGTphxbQtJ6
ZPChWiAJoXThKb4fNDuE8PoWMeW/p+j8seH5TzzL07sDLnBeHU4RnpEi5qQa/JV6qR6QopYy5rT5
yIwDvcy0P3O57JEi9rfgcDl1dx8bt01n61YXKGaA5CuUZ8nbgzwk3EZudhxpvuJkl1pDvrobwx96
CidsyY0e0AOSIEqb6H3dWbzvFKHnfkTEp/4na+2EWxASFpmlmAXwwxoKKXot693qb4xUiACOYEPv
Dr1de//jXOCiq5R+0tgMJe0yXgwInWc1/feUUUZxkOJF4Gfv1CH5Rjbjk1ZnOowCu3Fga5QdRvz7
yyuupioGhOmomqMWrZ3gvZxnpJwzZMNJH+THA9KUTnr5DCcLx0rlZBcrJ1utxWxFry/J92nzuHDe
w+4Oa/qgcmXanCMI0YHD0Q+z/aDqFqpUdY7CPSM/Zb7y93PqOeBaHS45gf3xlOvk+73cOP9RSWj8
wRx26XVtwYERcg7W4qnVK/f9Hvmm53qK0+evi75omw34rRTAez+x+15tEazSFJXxdEOaurJCfVNR
xwBWdgSnS3lNMtPucwXwHEUCWZ1mR6VnYOyBkBVU4efhkSCtZDz4wvB2OGm0vf2xFS6MAqBX1BwZ
SLFpL3sPuEKxkeFne2gt7xmcAloxf4TNPqmNXtDYKokST98nLGbtKJrsiuWteghtmU/3xhAof1rX
0x6f6HO9YCjKaDUbprtUx6i7uGYgOZ40FvxGEf86wAC300OpiF+/A1Pr7El7v/Jt8opdBJjDi7iQ
q7OhchVKytQrXaKp9Evq0xG1u6AQHgarC7vX4/Pxz4louJ4DrdtUzd/U6HmZBBSbrunR7RrHkNjr
lTuaG8WjBPuC+N93KC2ZwUCbxvfY4/L/i0kZZKrETq+TC8Wh409on2j4C8FQ93/9OHGlSTu5TKew
AbYsfmcK7h8flxx2MoDgt/Pl350weCHf4bt7xlRXHqO43MD7kJCkbrdmqhkS3uaxz7t2h/pnZIqM
yj0daio20gvKjL3v3TwFNNugfgFQpmF0k1YehM7DYHqJysulJ2eYj/atJv9tuGg5HEmY93ftpROL
eLajjuXxYUA7I5UkBWOAym4tbHhwmaUevcEOAMLvjN78/LlkVRHKL0dL/DTvB4EwxI5q0K9Kq+oe
dH4K8iCi5zqig2DuJ4UCjwTjHhEHtBX9qJZmncRL7ZZBAVV5NTJnncjzih/P7weHjIBqD/IVQKNM
WXKFJMKnJeJfMsRsGvwOuiEMfQxqoAVct9FYIgdsUbNDsEYyL8460koaPjivbgU+NMrFtHFH7cFY
RAOkk6BsTcpUD5xu9bTBlVTfRuvRQNTmpbNWNXxSRH8/cr/pSBDLYwzSLCw2778rjjqiVJqoZ6yY
dUbeS06zzhVvwIYwWXkmMpV29tp9zaYNEUpSGDpUbNDlXcFBxsbHe5Zyq+0ljtGVhLK+Jxk8ipio
cg2lTGhyTP/QPSA/KHfcULVlZqTkRpOO0iMwy1Dk3slg17ApHEgDMoAYMp0ll7tKGt+qzL4gzDGE
Vhts0hm39+UmHdAmMHBsnWzt0r2Q7gto5kspABVP+dYymiN7qxa4Mr6YDm0z9dfgD0aEm4JxJUSZ
bXiprVx8hnKutIMYVyWECa89ri8jAiuZVVtRv1V/JLNnpuLIABfHfrIDUpAIVFXFc2qHYtDyegji
5Hyfc5YRrneoVE254GL/kTqpRHnoeXMgXQCAKu6CoYvfnJnNGDjVi7ll8uCLuZabfPAdfK2ct4j9
z+vFb9QTJZJtFx8ine3BCwFDl+mtAS+DgbRKk9caHsRSjVZwEtywPCOO/60E/OyKeYkEWYeURUdX
L6v6n3F8guQF64+buEEdBE96r+1fwiY9SqfWtdYOdLCNmZs9wyIZoheOYDNah/Jo4+RA07RygIcR
X/vT9QgjfNRppW5gKWsi8LRnuctj7DWJTkDgYeVo/XCJrqk73cSWBocw+CuiAoOou9KUqVPfDedR
usv7OlTWvgLTnTNYqelMQJWuj98WTAZH+3qRfpSPQ6gnciPlX61PQ2hrOoIzUTLmYIwcvlxybSRe
WAuAMSfds6paQv44Ap3a1L/GYQBiEpOIzqT18jNeXsH1IiP19fnV0OAb3Yo+bydlpfFqA0/RCrGg
vw86VIVsVEPdCCogVvxGIaZX4Mxkyb/uY/z7izpd1kJw8cuDOwBF1XQODYlDZt/y/85O8+mLIrEq
pGoDuF5QO0lU8sawzTpgLjR95U0ZSTiJUB+b4SmN0rdMjEp4zyJVSEu+QhgbShNV4M7+k5gNEBIy
nifw4oE7B7GtGA98SRajxDXO5udLLQL4hhO2JmIT+NbJVOXt2DjuKjlG7i6ZDU77c4T5C9fuC9YH
YvsthJJtSs0RSjzDHDTZlLivLJ2ptJYPpL69t7Z64C4Y7H4S2AodJSvgYSemTyhSz4BxIXDhzBk8
Spy9KeiEk6lrkUcp50dBvzr8tu0WjWiw9Qh60v9KCm/qQ0BdAjdme4uSK4m9bhxIC4Y4EqpI3n+f
rRyfgsB1Vde9UWTh5gypHYoCezHxtHp7uvcvXMBbL7twpDGv/BO/Wu2A27AS6nq+tIpna3DGSOah
SNJyh5aIWP/Tj0e6daQouUMoXAGksswWxn2gvHNWtQPOHFtYd/mGSKKOPsiGjj3RsONHRB6xXYka
krPsWx0qo2eH7tmDFnlm/s0K3n100GaUwvUWeB50bt4RS/VYdVIRSu1CbBKTtPZdS1Xbi/Ra1Ico
bavUumMMxRzPKl/kG/YcBZe/sbYe/J38az5riL4cYAZnW4zTMJGPhLLAqabKg/SF5Jo6j66eyFy5
1gVJx20zid9knO0W0ud2w0oHUkPltjfl517Dhhbt78Eyzva94f5O23st9Mz49XvaeDXfPIXg8CMi
Pg4himEfr1uus0uGDiRqohzixnNqpuHXSP2LB1hz6hialN4luFd+0nZwE/dm1LyDUFzw8rJ5tVVc
XbgrxhL7yS/q62iVNrAbyGGiSlAeQHuAuM7VSM3351KQyWo6OxFGuQpXF+7H7pCRPxFMtIIMWrEk
MuTA4heVj1cZyjToqqv+j2isV/mMsqURCxN3kHP5maCLBJSVHDIcjDUsyj6zqmYcbRQ93p+iav8E
tbcV+sHBWQNB3SPIpzMZtHGhB7jpD6p/lNuK2GduIi3PzRu+cTdGy5wI3aaB7wKMsK+8zZ1eqKO9
6t+IEPUtqUu0SVNNRcboIkDa9A1KK4g1B/8UpAzvl9y3NZI/7iWK76Y8Owoc6XPmg1xRQTWcYXq8
3qxFTISd7VHrIm8ZiTMzYOO+dTelefSXqKZe1L0K0kGCgnjw+Km9cI5ill81grYBT/IbXd6I0eff
Gu+TrWjQ+mls+F1H9QhFqfKjr8AE/LGfiMjF4706fNDaJ/1KLQjE3zvX4p/dt7SjbIN07igtBsyX
7/fr4deXT6dptMG5umskcn/1RaSTtgEUwfJTiZvlWUcbzBtK+gnw7qaEnGSFUOf8E1q683rnUV2Y
i8WCQ+j0T+IClqBOG892dbNJvzJtjEt/9QzZLHplDSSD/lTsH/OpEK0IMNtkQn/kipTtpFtg4TIK
28g08uFXY764vA9S/BfjGnxVt/aIMTX2CBjIiEO8Q5Ycu6lhdeENNYdNVMPuNQrYZxCpILP7Os68
G6nNwI3lhFWLoa6OLolk+5oCORygCwWOCWzytEG2C2cz5+9v4GgXJ3I3tfo4/QaEU0Pu8H46G9RA
VmKNk1OpDDHHl7mWypjzBY27aHiOg1n57MUV9xX266nvjEY+/DS884zpdisA7rmsPpXeK5aKhOUI
Wko+fv+ftTIkNjYD/rohgl8LFa72ehZ7FoviWYgY5lL3+aS7x+95wPhGzclcTPUUAfxyTsSSp4kL
lF7KKKHXRF+gme+iS+ndsmbaspVnOfFfXiJ1X/GpOnAXAaXTcAnirKgGRkpyk+xhHPaF4JIY64ls
1IyE5/q1BtWIUPdXbi0GjY4M0r1Xuwkyo0IJ0fWgc5G6j1C5pMMFd0QObIIEc/Yii7qqXTDFOWV6
nkuQW1ei9ujnkKAgkm5OzMtspI0q/AcPzuGPr+LtCNmIN8TKzVR8kmvSTNgEjbpgcVcyv2ompnJF
ZHdP+rYmpZdgspz2ECiZDXdhgV2yJw6zmA7vuVgA7rT691OYa4UztdelaONejtyKpA9QuswH4EI7
hjwKEjpetRDdGdx96FjGb/1i4fdRqYvIu/mfFtFwn2+aa+ut8nfl8RVdG+j/ICAVuW02jvj7b6M4
bQal/u+xNKmvbgR57S9bx6nfty0ZRqlqomXr6VRrR2EL7uvZsNRba29ApJ1BXneFnrWgtKNsS5XB
uqpHa6xRJ+/yqT31egDUCtaiPZHQRyDFFurryLmes1mIfIj+vtJJHCzCoDTRnknd1ohC1xK4lW/u
2wJZ5+NrsWOfFGwngoYMMOzeGN5PFISiCnDV699nPwB8mEEhm7RFUE5zf2kgwmhBinf5ypvg9ngw
4PcARb9Ndz3yEOo81NcUeMbpRojj4U89n7BqaOAPRYidWZwJwbF5Q/h1ZpfFbUuNDE/vBYRtLmJJ
5skVpsDoW2Lv8i2qQYsfhWervadmTqujmeiLEOrar38VGxNx+EStym93nfNYU2RUupfk85M8fd7v
2Pk01y+IIphfeltlA8k75y5fRte7e6SGzKT0mWSZ+tcKFjqzgOsEShRqPLUPZ6PiETxPPZwKbS5Z
vHrnUoutbEZ8ypawIcafyeDpQO/OBjturZVMH/vC5XvQw8wmPbJkWrZPAHmx7PdxtH5cCa3KrlXE
r6jaRasqTdXR5i7m+vA1rZ8DtNmelfotUiIsVJpZ4+za8+eFgu9ECWMbUBeeY/HOym0NMzrvj8Md
dpDzSTrCbrR88TcDUqX+yi7b7Gu5oVNbDINRpiQXKMrDJ/ce+undpyinBy4OEq/N/zekfDmtyA6F
d2zy/IYOGHneoybJ582wESOMcwdAiMEh6rpc1z6++4g7nag/D/HEla12ckU4gg6z7Y8AJdsnST5I
OSEWViv4HKF8FjoZjrfcKQ/Xs6ctHFosm/YHoCZAyZxIg+Tb9ByZnP7hfZnByCmmp0HOB6xi7zw9
+OiwvswurjjIGTM8Kn9iMCS6JmiuYX1XBA3DK0VgsYOWFcKXHN2/N+fSiywzGKoqDzb4TWnhJhxA
JV0pZPt+lsewgkicLMMS1cCKwLb+3S+Wt7h8QZjI6IAtKE+b8YpnAItZxVAYBj14v3Hn55huIlH9
9aWovo5M+z3mQSIloz93eKAGTfuFMEICdoPTh2RKBGI64JY7A36aHvPIaOl8C8BN+yOJzgfOAHDG
FKzsE+xJJFC2vGmUAp2m0xuACn0j7XlwCTS/AURz4pbevCyKNmG3AujhYeeeixmXB2mgPfRYCJgv
klqznlUYgszdeJZeR+Ijr3wBj4sV2Yh6rofiEi6vgWMUN/MhuJcPgRBqgbGncpmCe9uQ+flIj/LH
8w0VJ8KJ8qelpL990wZyDW/8gL0RuLBlTo9TFdvmUJVMAweaF9tSzhngHV7boJaBgcqTYrYGsFHH
9SHXi/V2OI/4geC7eEV3jHGgNlRUrkMIGqpicdcOK8JWhjVUVCq5xzbNoJAEAjaAzK0upU/gw4mP
JMhkxOhgbfE4bgQK+erkPHYp47SL11/wNByUxzLKaT8yeNpD2FOW6vpff3o7zFyv1Jk3NlSD08fy
LRe0WtNEulAy8i9cN0Exu9KxtOKfwCzuQYqeUumJjsOqDbvwHIwsKDZOaa5M+CGVwXRMxcN3Gi/3
SeghGCRM/c4TT2H7nqlJ0Ps9CoJvqeUAWUqS2v0Qo28DuKgV75goJ7CWnIidEDUGvlbVU4DSj6xK
hA/txbI3gsb8Mh/PbeF4ajopMRDQIyANSCUbXnTwn9nL0i9rilaJtvo1GjbmP50Y31Jf/Zdz+zVw
kEQzNepzUBdgQ7GVc+wCWe3ayH7/GTh0urp4ayAcxcYkY/Wn80zCNNZ4OpGWFnXOMSk74F1rLDM6
BFFsaNEwAcJbD3ZGftmuKRnx6/TlUnwWqz2TPSXOf3HLOYNkTIMFqsJ9wUcncLXengdPxoE4GBaC
oDh559f2XwbUa4X21X7HYgqyckLNOmEHy6gFzbehh+u8aJpWYoXoVYCsaH1cjZG1iFBG83zAYFP4
QQza301MO5trz8oIeEzR7JhZcctGKkGhIf3ekR60fJcIY2KxEsIbm3Khu5NMrZUJgpwOMM2FjYqa
SEdswh541UVHEHer+Nte8OoSQWL9a/n4FLuMU50Y6J+cVcACd8dKrJNs0mg/z6q3wQDrpB5a81G4
Jgqt71AttMTZr5fB1sDEfSM5T0sJwkUpc1sdWERZr3TAIiVPL5ZzOZr9Scj21oV1wPHGcTF+b2tY
IqovGyrjPaQrwU5ROqro/PpyTunOv2LSN+C9QrkzDtzFZS9g/CYN5SwuBau2vHBnmNVN7j8MK6jk
FIFxCkcpLdaTUebtLxg6iytC91G7QtoRIWnKeCzVeVN++bTHLdgsatPInzwq/mjkiyQGZ5lu6Py/
ejgI+WPQXh0NdEbTozMVEUSdqsHMozNUKr4TuZDBVtxM5AgCyKX3fWtacKwb+LlYGA6LZYeW1i2x
a7t3d9rZMeWfKAMd7npdsRv6n54HZNq4z6C9hmOtN/Hxu+P1Nl892OsEQ1G33McAcOIWz/MI+jbb
oa/+MYibZxj8FC0IO22Momvg3nHhIXI3dS30lynDklwRJqErH05TK+QF228Cp2MU4i4EqE38Wqx1
uLdHMElE6eilI4eiLgMgeRUzNX6oUNg+N1HXtC7DMvqHjx3/r8qAM7zH7+sbiF3Vv657TcR2cCJJ
H1oo9FoHqAxCjuzkt6T9hMRQ0A6TlFV3fK9PZIrUnoA7VQVo9hPyGly/Fw2tmy10i8u/S1tD6BID
xE9S5WXXm0WFpj+V5l+7G+misxMC66jwsio5Oug5Bw1qGyBHPzrBM1HZsEzF5hZKgciPpg9z29ty
WDviewwiQAHMd2cixcqsD8X8cyo7zxDeGLSrBhX4xPu4nnwXoljJfNeA/IxUw5dBEZmXgP6xzc7U
hyc4pqp2ed/erT7IYa+b84F3hprK4NSUNvmVmHGLJtE5Zm04ukt0Z8zwXH50mCjBojKc1kXOjMW1
6ptaLRPwhrL0FTujMZRKhoFOLXfgGS6T/EbD5kHWEB/vL9PR0q2xoinjAj0re4zSsnnwyziz4jJ9
p5famZgau6YkZmOxnQaBWQM6epWCs59jcz8CadoZ4g3dpnoXSkKTyOXBTgcOTqASEjKtOqn1rk6P
0analzNFelQB5aNz8qZLgZcZ4GrbBNV6TKxGA9tlFYQkf/WhyrFncDILv1pGyCrbBInGk578cWxo
271tb5w9AM7Ev93mjqMf6rXBaAH758jkhlqw/6vImZqp0Cj6xg5ou2RzWdkuozUTiB8coK3LKNUz
tk3wVPlGxhCWKTrU2hR+teYpJ2skglA6SqPWz9XJ5gDTdE3sLC6VAz1icf9B0y2cMv2zAarb7Zeq
NoNoADGVAjdeeb/eHQ0eZAZlUqaB3qfANg1dy7b+llrVruUru8K5flcyu7hAfJdgXRir5F36rjru
HX4U04m0wh0hVKbdSM7r2bMzuk6C7A+1Wy/UVI5zQF/lQLMe+rcTy9uavzxttPq7RslE3bUJI0hb
ZJqrWhsneJEbGAUhw0il07dYgYL3VLmsfDS9wgPuFDgmhIOhnRMY5SnvQRDmV4O0HKqUbm2KlWb9
mD8NKNhNEMhiI3iWla/jXd5LYdWKbuEa1KAADa50dp42CJoKuWJZzzJ7ZRVorOflgIgjgDVlQfZP
X2UlET9mTs70rEtH/0NJRHmwpaMdPOEWKyiUkTwnuTK6kcgZnBuVIchLPJHmY/5WHYwu/mO54XTu
BAHuPe6MVg9gCvuOzfD09CKENnOTFe6wPRHlJaPs0c9Xw1ehRjgns+ZgOyPGd12cC7cP79HrX3iO
isr+fvb0TJfUfci6lKP+rU0bXqCeBWKV/0UHJO1HjnXRcGmjpVp8WJjpvmKFwAUUvy/TrrNmAWMQ
d5Dt3BsUx/phX+j+VEBEGlJ02yPredS+1xln9CupjoZn2Rv0BGPbpaNDU0/sSImsFO9KlQCHG9UH
FGt4xzOKUVIFVgErvyHxsMlk/C1ZdNOrZWKFBHWkgno0VTLZ/LoMMQMPGhGeBsiji6a7rpNO+wX6
dRqkwzKpZu/4bby7NmBYHxgFsiIXoTnOOPQ5jQUwUes2YeXJjBeK8Itm2FCTNzlsep3Ww7IgOF6p
kzSSOvPv01xEYyzPuXQuIaTkz4wqXK3ROhD81iv+GKbk2774JwKsRd85OhR5Gp8pfECueOdPvOyU
hxw+Qlrl0J8zqdLmsqIRIKhphs+rUr6tlkjtv+rbSQd9Nem5dootlBGlqoyQZd5hGbH/HcxcTUNy
KVNhyyzOTEVMYVH+jfP8ZreEik3ZHJYUA9TeeJ6Wmf1tOmiZ7XAL02C7yj9E54aEncQt6gOg9Tlu
LRsBxRkXNqZWeJVQCsJh+KSwfi8Nbkfw4KQOPnJjqBwJEhpnHWMqiA0rJjlqqfUKG8cx6hq8evFb
wNz3iZ75Rbn32phxqitI5lqm7L9Vy40LRgtWjBIysCO676k6dKx3K1g2pcKeLPMx8eObQRNJB//K
5SoKlAuFb2LaC2HokPhTrpYKKy1rbRWx0lU5Jb9C3VBlMk7g+iMXFYOJ5X9QEhxEpTZH+5Ik2UJd
1gT+Vfplu0zC7ZbqQZ47SWci5WtEr/npbBGB7QT7ss8Nbjc6GonblYZBmyOl54nY3c9E0OkSPaiM
1Na41xS71sqNa2f/aCEM+6USmUDXfKEKUwnt+yxaHGAMYDWUkfg7FUuOzi+lZWiLRURVoUPTdfCe
ZvfwM7pzTYmUOkZDw7OAroytlTo3A97OjI9Hea1rMsw4jEA/VIqJ6JXWbHBlWG85g6DOSqULv2gE
D7+VGOSVU37v+VTPQ7/QoYJDfR72dS4qyfEOHJbK0ADdpm/SzqIZuNbgwStpKnCSNoghkv+1a3uB
mMyOjMFqEhtryfqv4UJeMr74VmjYiTBaw0FM6fCgJn5H2Lz2w8jiXcaHVj4Gi2ahBKfacMdUrxcH
ntd4wq0dTcn0jKD0iR4SKax2ozqhsslS1ETXvaY6RJjLFCafqMUsWrgll227g1TRKIYbR+UR5w7t
Y2BVdAtWPeI69wXOhtC/mAwBJJdQNscBif+icxU8UtzWcvQaxmuV+PGU6o6UAa0UPuzgmVoYr0Lp
G94oFvGAjU2ARpvLOfy3chnVuoP0qYiDdnOgUxCqao2TJNNkb1C9H5WmUSkqEHQpE6ts1M2hsHhL
1PVUm5iclp2SlEXqGvEpVShjRYcRHvAwb7cszq2Titrr9UUi/vySgC987y3RSDuio0Io0yswYB0t
6JCOCGQV7EDGzjgn3p1B0UXIdmYT+rYEH3AK5pOiGrqwPkLSJkoxdlmEwe1S2qFeOkJr9zjqwuwE
8kpWrU9bsQh8WnLhtLH1oK02hqNq20bTw2iYUfhvQRUrcUqJ4Q3xQSFBDRpsykwSNEFPd+rkICR+
dMS9YKYISz94ZgoB03XxeW9JYqz3cYLRbT9WBjUVsaMAEmqzHSl/qOl12Re9IAhjpBTwpIrJ6yaJ
7vbzJ+NkoZM9T9FPIUWSeIbHTAzxCBjYWGHokfgQ/QTPRdDYKqgU9N0HRdbX6rhKca/iKKlDd9Ee
e/cA9AeieokhVR8PwVqsG6JwSHqB+eMIoEK23GEdQItklwZy4tMWFvpd5e9bdbckNabk5Y6x7Avv
B3er7Jy/nIzh07H8DcATYSDpNDjoaJk909UIxti9i1JGqwDh4g2h3sgLKDpXAh4dQKlWO/23RwE3
6LS6CxJiKLvhV0VvdS22BzXla/sfvwmlBmoD398f3rbJPJSlKrfjx8o/f6QppEmoHqFw6OqYcOVi
C+ORrE0CezG7kqO+Jr7KRQJT1sl3vGM+Sr+0l1Z5msOaRqbtfDqyAsEG6yzTw67R2+JQMxJY0iTK
AxkxPWDE4scbaMIcpY72kzIxo8iOcP7LwGx4wjeyyN0InmItNDJ17mNBEoc74D9kLKz/p0NwC6FS
31bqU5LuudaHd6+9ooq9CISeeyFUwJAsK+3XfqNeq3O1PGQsBSa6UZ/k5GyBiGA8xopIlKcJ2EmQ
BHDLVGY75obnslXrLWWWseHoNsnwRbpnzFfLwG5pyyjVgXIDdri+VqV4z1lxp8YW6/BcewSdhqgc
gOI0rQK6NHmG69tb2pD7UvzabY0wLMTxJ+uTPIcqBNA+aQMZuLwOcIxor9nFVOS94nnwGF8sSa5c
TF46dhUZn1sPkHIKh3nv8RHqk+VRBo6c6ckwFNZ8PxaQTlh6ASzzlwVb1/dhfmIMQoUYHR73pRns
8NjvYdgPdLHymcqK7imR5EK4cJzGtLeflaSoGcu16tJ4iamav+3P4yAm09Akgj12PpwJ3lrNth36
BW65tHE/+lWwPXY6MCQ7uu/M9FtxGDDQIcxVpP4HHHhf+6wfvDofEoujtiKp9wBdLL7Lj2CROp94
aDgFWosghwakZCdz9j09PZKPE8b7N+etf03wSIFhNFBgJiFlvvmQcAxdxWWm3DVVn0ZmArp0Uq3r
f6Qp99D6nBVKys/X3u5TPwbpHv3kvQXvW/W8bUGBkefWt6P1669JjUsOoMBLUglgZXXJiUGO0IC3
m3WQuTzWTXeH0q1lGhK95FjrVER27YSYLOMrYUu2hPgaKLzxqHSn0A5xAab2tmU4pYCKWxiQwmf2
Nye5scKk92I0r+5c6EPOGP0MbNGEiZ9vO1Kr5PjVYblxhLXFqbjIawqdib9Onmc/hDFaEPkfRr6s
7/Ag9jYvpsxTYJbQbeGSWJz2BzbTzFKhAkHyyWHjx+rnRzK888GVLwG70P7kpK3m7COuT4IibPBA
g0NK/p1FlDNyT/O8SXLaqaHkkU+WnQf5hG9PB2mpzs7TFhIi+dyFC3LaCxVT5bS5WXCcXFBRUl0N
+iybILuYZDwhkJHOfxKS5k/a9rEQ8Yv3ULvYNRSwx8zV7S2HokGdcGKHL80ktb1LwFMji3F0McQp
CrQ4UJ43xt8NFR150yvKgdqDZ9iM8fGQgJv7CcV+W7qUdSgZNx8H8oX89ky4ZJhBlaeX0f9xoThs
KCWf7mJOLRUxnMlIQuVKnqtD5PRqvsvYxMogFe2Ht3Ml1DyOI2RmzKABxIlOdmSCbDlNbUsYIjmn
lm6djf2Dxq3y+H6yuKpVy0oV5E+4FpKdumpLJV4fflHDlKrc4SDKYlTBjPzTTXD42Y2umC8iHdgU
V0qJ3VMN3G8g8ZblXC/4s8FG9xFjBZXR0WX81RKjQMapmSdMw1AAdwVOt1Js3T+07D5lx09WiU0Y
l5DI64pnYtHXVxaR8IxtLe2w3C2rdOgVpCGiDGCW3FdkA9+iIio5snR1LEmKnXFM4pqoB5lN1doB
ozlXaHQBWNBQX2mMu7Gs28EdagsVL80Hh7XrujTGWRklVSpNDs7AxwnZ/t7GoLF/Gcs+j8065i2T
+9avDUWlWVJlb0XA/L9vn43CwzjMyIupP6jiHdgtF+Bb7bOeG+VvBYhIuembBaIrHxZC+EsCGKTf
0tA5Iv35iU33m7gKOAT9epXTWBHhbQDklCpFskUT29D6mYGTqNfuKsfGinkBju0nE8D5RusUjSsR
AvVW204TYB9ayPGXOCC6FuOCteTG2FCeANFx5f8gptZRBdwzkBv8s0UYtDhkoHUm2NRjU6zvIzRt
ocuOxstkqkFj4i/bzyLlWVa9h8Gn/LUmJp3PiDsW3qnzazgx08k+AV2PJ2gxmp/YM1HjkxTZHTCM
JhgOXt69nqAB2pOZAjAbvApedN+mBwIobl4WlFKBNCr/mbOb+fmNai8diqB0UP7TsXs9rONn9GEG
tbYzjkIZMI8Sh0yxpTVr95cp5nEFbwCP7It372r/jwVWG4TyvAgc0FYEll2Kr2abHLzZtlN69iBv
ZS9aXpl54sCMyMc4Y806v5Bpj2l20qYfovUleaZq+Zzbi1doG2XGfkwfA34y2PRkLYt+/A4uv8oJ
uGN0O5YlVgIL7b2Dk6mdiMD2MjkXrFK8soryJApaJdou0DsRpttE2sEUtw9racImzAGks6F7r97q
8VI18HeKc/XVU9t6T7a46W4ccdse0E045O34/gscOsvDkN2mbmFT4ECLJS7LW8N877HYmT4KGhjp
3ioCfZ+QBv3AK6+TSdbj82o8N96G+L6auSchPurTrzVeFDZYJR/iTD4jDZ5V7hGD9EiviuHyRs9e
2Vmsrh2uHH4Bng26OdPoPXa/SECNRWn3wVFVPqOg1JWldDDybcsOGb4B8mXl0LObK1yGWUaidqv8
OvwenQQ7JeG0TlPNperqDRD0/761ifCV/0F7eXT0N5JP8m953cSOcJY/un+YZ+5WunFhQDtrCIE6
KmxTWCoayVIKPNRK9ZjzBMe50IsEssK91Sm6NavckFCCfG/yE4DQVDcrp0Bl50PIAmIzWmAz35iE
HJlq34mk15YoxwrK9DO5IBogNEOruUMhceZgqjIQocRPLVRG4sBRA8VxujXJQOzZztXSR4qpkYeo
tcXc5fXSS5rf3vTglDRn8/VGRuyS1b27ZSf/hxxYiqmlTI6Ju+v83jOEB+k4FsnSjQz68TUYP8To
yCxIAEn7UoHDMxUKu26yUrongFBJOj0T3w8BKOx8tVOynZ4QLPtsmYmD0Gcqg0XP5yJ5GxkUC72W
UMyImqWHPB5NA/X8XrY/tVBUVoWrQ8VNGmEU6V3Ow5334qpTGbDIg0M+sfOFy8Qq3WpGTRHsweii
NrsanHXLZ/n83lYvVdme59rtN9aqhtO7J6FhAqG0fmceY0ImVjrMqjStHoQSkDkd7qWgLU0HLzxT
5j+Wy70F8ycmwUMwdYXb39JFMOeD4w/4uDYQYZCmP0tpTVjukXlIWFpS1yR7sYJ4CnLBKp7QMDAN
ZsqHMS9sTnLoV5Rae7e6mFsHnqmP5wrM+isR4HuWjoH0hUZqAZH060THSphjwsMF4pqWRvCAhEl7
TOweBG2MsibZu6mE8QyOOpF/Pwh6P2ZZNHm6L8m3NQbPI4YyVL24NuCe1zHREdEFZKwcVhi0gysQ
ShsHQrO6nk+rro4lMXVqOQ3202ndrN0rwt4PlxUDzLb/UKCVxu7i4EKp3mytF2pR6fu5oPWdhUbA
Yi+/1H1JZ0rhrTkcjTAHZs3uW/qDUCWaMCeVLclK/qFY41a3zZvxBapqr8PQo+/3WKVyX2j+hiXX
rKI5561t+yemkeu8JCm/6Cnk+iEaacz3DvnA4gxxYJRcBdpatY7rakst2Y++8V7ZtsJVn4PR5cOh
gBhlWT1+36M/qlC0UayvlXN3qg2uYcRZXLkzk7K0ySuMzm2NT6njojH0/WE8RtoVaJjpUaVNNf34
yEDAYLAMbBkxT0rcpZ7GWa/ULo5tokV6ky9BADPVBdRdMZjTTG9vuwXaOccDrxHNMwmEfTr22vFx
VTMuzpb8ZWJMHvwPWGA4E62vw+lthw1/8PzQcCqEky6sSOlTBF19RlLbDFokBwjw1K4SlMP6e0aO
F8FhhQjTxA6sScd9T7etKsd7twdzvE0ZL4Sf+0J4KBp9hAx+Q7/IJ2HH+gwKaSTd5KQonR0Cr0bu
PflfAbDDRMXQE7VFIqIhjPNrQ9ejPNqRt0y6bA13MLXhXORaBmrq3hZWdTSepHP79z42Upl8uXHF
i5JBlEjMeHDDhpODyzR0SiwMXCjSuUPZvZn2TI61/EytHffXlwQ1Lbo+GQTD+Gue6RANoiNIdc6D
8VWrB2fmenOOJoVbsuuYMmSQZI74gAXdTqnpfvIJpgSvpokj7SqAZPHw0Yd1Ecc=
`protect end_protected
