`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pNwDVGRAcKAZWXZIVTSVW9M1ZHH/k+FUn+iq6Onu6ngQhshzAzqAa4tbbgIVmPbaESnrWt03UH19
Sl7ZVQ2GQw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ejMIOdhrd43dK+qlMfl3BrmT8r8Ofj1N5k8xM+KRVLdKfj4YNx+3v7VEeSdPdHTdZtJwpkYEsj5B
iZfwaiYxC/AFVYgEvU2X5g4pr/rhFEUapZN96pKM1UEZcfovT8uCiOnqsWSET267UkqISGSqK60A
Unm6OfPPUxFWWzZ/wM4=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
C7xDAtdOGS+x0pC5MvlIJkcPK4i0oGA0kMJ/+UF0keUE9NSNYygaftWplgcQ8v1d5tDJA/zdsozh
AI3WFfsP/IlDVCXHo2H55+352yrD4+JbJW5Yh8K+CNHh5AA02rKx/dqpqqQ9BOgnqxyHygK5yFbz
12gpQuU9InGczqSjKkM=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Hf/oJoZuhJn2JdM1KQwKs3D3/2n27f+Lr4bRGbHxUvbKNxsuTv4b6ua9w2KjUkPpUIcy/t1MPFHY
JTEYtnWI9NkjCaOyNyOP2JgjAXDzqfxi7xKrrSu3KXWrY56gCCMi61G8AAZgN/V33joBq6PTVNyq
7Mee65ZX8jK0G9mlHOz9JtXq1Wl/0PMRM9YXwQH3PiGDzHoFgL8411yI5aDOxRMocO5r40fJRS7b
eKyUJwccE+QFLatd69NV9BTlk1T6BaimywA+u3E5H6gL2ddkCGwscVE8iqAbzk8z5ejpXz7baJCh
rPo0L1Ou/QpdbJlDQh+skh4hwcrR8wAvbbcnsw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DOXSTl+SqsA5OmzNKMoDRUxg5AkLQknSJyjPcJhpcAmhq1YF9vluej7Lf0OXP2ipzNYN+CB1lR55
kjUbEjffGhEzPZbz0x//NQyzJ/CbqkYQqKu2Qdf8RVdJdtix8SWELlLXv0ZQoTbe9R4jQJe0zMqt
ficm5RI2Ny77ZcDDFvX9VBwfpjqCNzJmU/L2ycr1ApYbYHOiMsqQFUXWxgvriOnsjxJsVwcqYocx
B+6qg6CYRrweUNl+HqRBQTQ2GkMf+kWC/TqCKEOBReGCHo6OQ7aRE5VoKIMBsoNFttQPwzuQrYe0
uZRSC1delNby7cGHCiDFPlvq6h2lLh09Kl9cgg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HDprZpKLv+h17ED7/4M8e0Xlm6OvRBeA7PvUiiVfDDdm/2f+/DQ7RZ5r08EPY1GsewAdyDjmcjJq
lptnuj3ZeiPGwvlEqD6FZGJQuLfNDcfSNRXuna9rH/FAkkx1dTqXeUKRautfGYDCsNccrQqdpzNv
fD7zTziz0b9Ka82UVuVFgJeIZTpXXuy5R4rD8sG3SP9aRBlgTsoiHW3LIptS5sFez72xKEsi+xTV
DOBpPUJImVMZwIS4k+vlXvYqNvhqH87wNtag7/umeO12UrigxoMSCpP2LlSHCOS0Ki5iuCLNdtii
jLCCsf2yge9frWoWPDquMdgaWJo0D726Rc1CWw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99632)
`protect data_block
Xxa4gBk4Vn3/ClHe03IS9rs5itfDJjv1EF7jMmaDW7aTrsHp6ODOgTfCGPcly8Tzn/AVmH8hELkO
1yCoFUeZUPrTz7O81ki+ckkhnL2B2XhG2/y6V+64enGC3Wjv0a+hWDeTmsAvvEs5HBkEgS2IQ5f0
UBNjAq1Mis/WXS1PXA/8dVbIqAQE+A5vBma//p7S705J2sItxpm9HGG/eKXCAqrpAr+LPRqLC6je
DPdKMjH8k3SkjZE/Axou3rMzgUlj4DYwSxBdumzi85gEMmqPlUcT1qWc3/UeGK2xrNvVtAYtnEMY
O2JmvJU7OHCrQ0ced2fVxwSsrUqsigfWul44GpY4/iiXZBXFTmCLI/SOPXhFkPaiPHOz+4pbTb+R
KzEu0/X0LgFXMRx7o+faeSPkQwzjrlmn4UYyeyxo7kkkvyAGYYcOOTY6tD7ZRysX8Zj7UI5TplTw
AwMyAdbGHG8Mi2vaq3/ZZ9J4pC0ZqpAmwA6tF9RqynDf0QL5C0tu0FHNAf83+qHvhdxiFZqpFfeh
pQhRXGCugAU04pFbJ4muuYapp/d0WvkbHxQOB9Q7IfjoPd12xcJpq7HJw2egvTOaGjMx04YF0rYM
pxurWn7DYMeuU7I1ZXMgYqeCwYzAKPpXjVN/ddg9D+occuDsaCF6WDwui1PqPOZ0A11hfoHxYdzC
f8dXSTOabdLTWhOVLDjk7CczNBAom+CtJAYsp8dW8j5FgRyItc2AtSSSum5QAAcQJs1h0udS2U/6
gHCNRv00Uuo7Eq7A3hAzaoWxeg7PGXw4cJtFw9XOE9wwPOArKqxxQLKtQxlqOMdOfKc9KDspYCyq
5nJ5GCxRSHTXA1Od1CDqujzoZM0Kh5xxmIkUcvj5my7yo0z5Pe6BraGzlD0/IGTDtmN6PeMSkVHr
SEq9m4t49jM82JLwa5EDlqAtbvtBuBy5MaGSCLso+kNrjrC94CWHWE871e2naR5K4l+H+uoRI0Hr
3/NikP+rds9NJhHKtVDk9rvizUuuE2yjtIKZgvYKC10QtAB1dvrV3jJOfKP/UGkV9z6l63D2NgnC
kTo7IlRozhmWiH484MmxH5WBqGYAJpaVG7ZAy4fAzCng22HlF68VhdilMg6SGyDEGEQRUAFFdP4W
bVW4avJp1545UqbnIf1eOTl9UxoIgYDM3KBq4KENnF4vm9WFtvkvz0oMk+jKVuTS5i50AOGnGX0y
COpRvxIaYkuvyf1myFY9BQbkSCHcyu+PHaSIra+g0tTeKlDUemTcA9hvtn69rOeRdl0WPMUZPh0O
Fqx68wldYGdUc2LV3ewGj7r9M7zC66uUc9Glqcmrwtn8MaX0OldJrnDSEUIUvdoPmG94PWTQ9/P9
KtLnsfUGVe42xKmhXwMG2c3U/8/YSwl/RAY50n/B2qrTk5jcmJGPpO/qCrq6Em4P3erjgzrqbhOX
XF5pAOozHlY/oplRI9Kzx+vUDpuRe/aiNVvzUxzL0i8TAgqnx/OqJOCdGncb/pGYcu57wF9ni4XP
SzIe8uDR6GF7/6LRU4Hm/KkfqRszVT4oXKw25I3gp5ktD6gFOQVM2pfciKDl/0FctXurHZrfmGql
4SMWk4cL5neXuaOFgP9jI0JH1LmToFE2/RlGoM8xpQDLKjzV7GE7IrmYbPLFmUul1Sl5et7R0OaH
Ogb3LdRU96oSGrWaOuAYJd6r5Vq1pViETzqCt/p1GavpoEEhB+ZzRB/FL3BxbjD1B1dlu1BJwfNr
Wm9N6RGZNj2Ca3FJFU1ZDpvZj8wrsUig+gMT4MFsGZimO7ZMhupvzTdmtZo3L+OVfIs9bv4odU6X
5JDdnsHKdIc/xNkuaXn5GHYSw/vGvtb5VpM3+TcXn/IBMV4qk47SI2iFQHEFpW7ybKL2wgTs9/UD
DdaxUeEa6s7Zn8By9SHiqafXPYdqNe4O/S0Tb1+Wf6YA3OSoGQ499obprc/Sp/q7b82ZE6le9+yb
6GgWkXPnw9ww7ifP2C5HrJtggrxwd03/GLrtmu5C4VsFIXN6zVMTlKEMFIFAG6lZWYU3UrRDYFL7
nvjnaHWkR1bzSf9EyD8ggrHFCCS8kq2jICr0zSlDdTmkKNC7h57WR6+7NLtjtsUDYFzmgbhGJQDJ
qDnGKkcFufWdERMVl68jg6C2MmAwOP7vaP8ZWNNB8SnQwoGFLZGdLS2UGBAaIBZb+xHneBbPkly3
qf7H+Gt7okX5RESZHlQWzza8x57S6ESr5WUFQE0H/4DGz+sq6GarIzLOdlZKSPceQc09Mta9Upde
OKhI/DTChZrbwPknM7Z9geCCkBkRWuLqYpCqx07iKB/FhNeq0a9NJ7FHNLFjeLGljO7nCvpzDvUv
oC3lPwHR9JuIEqr+4BIyml2y5ZWv0GCDWKNihCcHTkHKKgRDvuNxwBKpv2MLmjXM9yTrABsGeyK3
cOJnGqP9kvVVp+WOhmyq/rXxxsyDGVwIc60ezjA5czv49WwEXEt7g9MQ+I1CGZodD075pG8Ygi+0
zqLYa3u6lilcp6H29r3ytF0Y2yHoYEMaC6U0zTd/ZaBq2iEmHTLYKaSdhHpoM5mHxBxaK2tyc5uk
ePlfLHWgLylEhNIul3VrN2TyPNJ9DQgOdbjiDJbHRlnAeSJo5Rwr3kxZQ/FrcFX8+TEvlOMHLMVm
C/XbpVy/YFmwi2dsz59kOuT4fEAoEriCy72jbVcyQhENLldxuBv6JPxZlD71w0gaacDsbUFoLLY1
oFlayKhrRagusJk9H0rLCirvYFYVc1wEQThgDDQCHuWIz2bAxaYFBlj77uIiVSMc/Rll8462goJt
qEijl3DUCDsU++ttWdCxHM/vlqKxTvrj0zUwJ7xfyad2v00YthammglpV6iPqLUr2FLSZfmI9ClZ
vUOzOXRZ+QQTG/DdjH8Iw98u4/Qc/S1ThF0Wm5QGnW2iZg6Xdvx3LwJJQHnfZ2ixocRjc1ne8qr5
FtrKssoYQNxb5Q8PaQWcL327/DjIVsBwCf0aYlpwB60boD8LDuaIdkUgZD5X4tbk892xHz7O3rYs
NJTx8WdW/coxJSWMnKsp7tqsU+HX9vTQN3MOQw/aPwo4bVPxFVXWdMgGlnhqoyZIo1zJz3QP69v7
kYgIuAyiQrh8SaPj7BQqV74sEcZenbKhPl3df6Pev6vqWprywYWiG7MiM/BLSFkscf742mO/dIqi
8emVsR8huCE7quY3LcAXn88Agvk6cTu8DBy0xi79q/zkt6jmD7oo1knkeIlN1TSmp64atfboBugT
XkB6gs8OIU/jQuC8pgjoqMNgcg6c8bLzyMGqL7RT0s+uqNQGCyWT+rkxKGklnRJKTJBq0F7aUr+U
IWR7Aoen+jmcPck7n0QgfWpnVRincZ1XKNtwOHXNRXoeYfCQIOq0O9YAAS9ouz2P5F6ZZvhhaI3y
e2yNq/FAWLwdoaObW1A/mSyER8bcslEfVxeetVJz4JJ1zdgyE8ZI4++cdp6KcyrC2F3LdMfXiI/A
IjnSN6ldO+YO0UDUHA+jtZWddiepJ+tNVloMV5uDlIiFKUfkTnLvcB7Wb0Zy3m2AAdSR8YPh6J/W
bMrkBmCro+lktp6xxW5VhcxPQjzeI0pd19FdBuYEpUXXqpeluxVZ35S+bNDJSW7hTg7F6HaP00lc
KS569y7IOjRdjOtJUmeK/yW8IzDrUaWjiVMMTpU1uUbGvKBy/UlCER2ONnFWWULJ4voOu4F/XUJr
lb8xtPXrP4/RwOs8DYMH6oRjS3FoLRBv1nauc6g1zJxBOv59dYJAaLidgph5rR4u+v8nOqsqHPR+
PFGgHI8wQAOxJhJR2Tj80/1+td+0l7+qR+aMgIQJQMaHzY+ZmpTS7QCGRSXdAK2Hw0nTeeJYu7CJ
Zrg+39yVH34XSnFxpV4KeAtotlw5zra25aFYw2dVga2oa0cTZPfPj1lGyZD2UZnnDjrvoOhXqiym
YAe+qbQT3Am2Cjs2W6V+OcCp3+9iKYpH4Pslb50cY1rgK2ws/KGjSmXnFxe/PN4intbmfBj8EwHw
6ZjGrfSU88fGUfGg22aaZGk4XwbWGzjKpeqp+t5w8ipWz25mlHCLZB++rVZ5QyQHDtIHtHsvrPon
Dn3vqTDiWUysE9eNWSU9dHnTcxuoB/4nhoH8mZhwsI/9bMoYyFHZLVQjn66AqyjYyOlQLEVwZ1Gl
4GXtVUBqzldQ6NVG8NwC5TvZeb25bvGEJ99+W5h8E65Kt8WPy8LA4N0z4emN+SsyWo2A0WLimDYt
FvRCUq+uu8Ub34SN6YNZ5Zohds/iC4BQ2gOd8tnsENUVdI3jJlEcId3D38cFs7jqg3KsRWnUXkk+
JlrxwFmB4a97DWLff6AC5AeCTrgLOMfAZENgH1PAHMPUXuNSp5tbhre6SK0hRIDSkf1XSjESffuX
tcENQG+FRj9ItFp3Ov1VNmruXjOtcyGW+fyl1SNo7LhHyjfQ63ODKeOvSW/bMH90AGVrlrhjbtyo
jDfTElT3qxN7Ta/m3iXMxEH+xsdSKId1Vq4MYSnEzi3BSv0vPZD2vakdFafBoAIC8ANWRcu0ZmLS
5aO6Q82PcvXIP/eyH0BIgy5xe7SEUcf41kkMeowdozgOJT95hI5MiEjo7VcUu6aSZFWvgMIcAKaV
47aRelaBUymgmowF9vv/es/HIm1AjjfI6VMbdarjHflhGhKCzdrD7zxOHsaouCQ1dx5I+JILk8z8
dm8oSBJlx7xf7QP31OOBCi2N5bXdoB+RBJGkPbrHHEGy3OgikaWX6NNk2aFPAABWTUYIuvi+ELZf
iu6KU0K1UZ/TZN25Zkx2FW7gwRGClHR1+3YbBl2TPwSvpviloH7g89yHdWKRR4qqxlqbWVDvbWkp
KNYE0l6LcUvOVjnQ0BiEQ0sXDFym4nTsWIVJZF6uc0wVXFoADTG+kD6hTWPcIQKaOmNTBZxInyAT
TrOEqp/GV0SKX2Vql741xYFoB5+qMMvdSkR+NnWUMFPfVUWUO4MmV8UpqSNAXGDpT+dSot8+JvWF
zSNG2qMQ40KuGNg5BzxZKF3B2x7GbDC/NP58HQWBFuCN+eGULGq650X6kFMOIrFW34/qOEXAG9HA
CficI3hOZd572NJk57OvGSaxCRUBZXgAHZKnmhNC5rqzH30Q3bCJYUSFJgrbmFEZ/JpdaCcNSJZj
S+CWUIwsKD+rtN6YrUV3sb/+lZOQUNDgK8sxrl7hxkLb7bYDIx3k4JOpNOecosSQ8SB79bR1Qwhp
vSCuai1+DCHssRgNJOqD5TdEpAqV/B+J+tq/EQH4xoHQI6vsxLU97Qr5t9CQhV3qwtN/CxcfbzJ3
L/Axuw7y15CFaqtjK3y/DXI3H4xh5hR49pDsaSrwG5ORkCoYuSDtcK0du7It499KB2kzLukoX/dX
itI7aAM26lbi0KBh2/S+7ulmTJyiSB2jRXgLk2wsVmy4iy4UQiHC88ds9KUL6aPU+fpAyTktFaKu
46mPMN2UlGzZ3JMMcC+Vm97C9qqa2eI4Drtd4ZJQ7haHNzbFDyJ0faLDkKTPkJA8GGlVge816et4
f6hXPYcx2gsOkHX7AiVZCYmmd1SZpiP4lT5XzNOPAEU7Q7wtq/+IVwtmUYDO7QW8Fam9hVhXv82+
VGYCuNl9MyX9xcLpmey+ARjIFwN0N4wuvWmeYhSQ8TxChFKGjbtEYz1tchfQ7SQ7oKCjvPHBMIip
+4Do59IbKT2HmQ9GoC0S6xJqXb0cssIw075J7soXUi95uBQAnPyIZGlT68ffry0emWlu5uJV3qzr
4J2GJiNfEfNwH+xiiZAEqDG/85RRjCljb2Bg1TDVf+mAPqqWSDyFriNUh5+NXljOzkfXzKc+Kc/D
5PWovyygsovWCVwjhwtzUmrP/kvllk1Y16oItbCIJbPRL0APByI1U0eVJtLNS0ITuHAxbbU7UGqF
w3Mj9qwTy340m3TKhjnElmTtDx9zH4KD++e2kN/Gmbs8+w6Xr+HE8CYsnIzsYLSyGIGQxEwsszAA
LN5cb7SkLDzRJ1UjAdU7abQTqXPTGjsmhM+tierk5YbZ8CohFZOa/GVWml2H7ApcnwsWruV2M1CC
ljI1pqddi2L95vQ2nWLJHr9kTIgsThI7GXh+lYoTzqP9s6Rmpa6jSvxoVl7ZOz7PGxYRiCXag0fc
KTm5ecPkg6uYhVe0GrOnQi5iwIskoFVakNlAKPmHZkAPkL8h9DAqHbjBBXQSd47N3VMAxRtbSPrR
o4MkQTvUKsa62P5wyCh9mpsg/OWOF3hcxmxlWYd+A4Eor6tR9A4qMMT8zB2JE2fnYHJ81hl6tqGq
AMDRtLX2OfflEuzRBF52FIw1UaRoibj4KOM/vIm+HpLH0c6rlSPoyxNkYS8S9+KpJG/Y9RLH0loe
ayH8mDdNMgGKdSMuER7tdldD/Q78vtLjzdpWQHrC8ChLsgsCPic0TEAtqHrAz7kG1mn1zmAu/y0y
Vwh60zCSw3YFkR4sCBqTZoAQBZ31/vwW959Ub6xitM1nNQwfRcK48r0q+AVI0/imHZZPtzq5s8gi
EVXahli9l+evk1GX0TnnOddE7Y1qU9KPt4BF0ww9gEf9LvybfrU+D6r+Vd1pi6vDEZgtwfYEZGiJ
fk0xZQ6UmAMFmdDUx7NMPt8lvTorNXJ7i35BcbqxzGuy8FlraWN+4+MutQ7E/sX46JiQ3D7H8o4F
FGEZ20v4ujEtAYXPU0MOwfM8t0bwmLBrgSuEXzS4LvkS+yvUpqsRg5+1qeslo0oVmt3fqUzQpOq2
Q2djTToRBOx9fYn8QfEuKPSpPToFB/nCu/JT13EHNXqmY2QyPgkB1FvmKi93Dych6ASy2vFxso9C
I7parbuyaQOVN370FohfdyLhtO+7BFMYkLv3QIeF4EfRMgC4t3Br+FDu5zJ4VCLygs8nl/HUb1G6
cXqju5FCNUGW8ro/XEzfT37nd8ng+ae/Ter6Y985+YWXVhSPhj5F0J8AynbttehFtKgIBTFWbKUV
ED5AlIJldeJo/OpfR2zE4cO8aeIsWyb5rEzmm2kdTnuc8u8I8gNVXntFe5HCzbGTNzeodXHAnPmE
YaakwL651krdoSSqt79dV+UdV5G9nkaVdhuJEDIS8Vi/ZpabF6EizJucvVb4nHoCmKyaGsOIulwE
aeDvT3wK6xWUqydRfCjyBWEkce/HmJcxhMAIpDct2KeS2+p5WZ1iSyp+e0Ct2BET1XUpDlcYtuPd
lDwnKKh/OLsZVt3oRuk4Wa2qJD5lXwf9LFz8QhLIn1+q3Bud54jbjh52Oq6OZHrcXhFs1ln+J9at
2aw0K3vxwqsGI9NP9vRVZoZrgW1eTBDaKSXjgxUr8yS8s7MkQMLVGB1mGAxPKCRMMwZBVZ2HaCm2
5yjpZ9KIgjHSQaNzXxU4rMH3cAemmS1XcSoMshkUTZWXA1CptfTTnajvAXyimkLbiVIeLFMbT6ol
swqALMpPVmg6txLIjTMKkwWB7e62um8X7nVmU7B+ojZ5LdUcamQ7QbpB2ViuBmjO+jCPUVxpRpZY
L0wWsxKIQSUfHWu8XuJUyWBAQ1iNtPNQ0bK7mDsspAdCjMA7aOvz0fZNvxMuaCsdsZNCrhFtRTId
St51CaIif22frUObvy1d6pFF3znTW1djkVQ4WCX9i+kdl+D8KUXfJmSM/nFFDIu6V/sX8hu165Nf
+huHKI3g42JIQjhFzh8QBzZsUw1UBL8bCnPwEcvC/6OII722wFLBtCaQQ6LJzttffzkptMfAWkvU
GjqynmjuHLcxL4grLkBCyaKACa0cDln+Cjt/aPyhodr5M8tS6syvOZ0L3zOjXvySTsWXVeu0I6ek
tecQpjIg7tH3C1MMoYDp/51akw0XeQxPCnKNnryuOvzef+qt+EBhY0cDio4C6drJKKpJN02lknxZ
IApBlCtbyxsdSFz01at2WR+qE2AdjnjpSiuih7mr9Sm7gLj2GLgzD7FfALaCLmIDRmIyifYsj7OG
g+30aJ0sHx0d6uEKg/bux58qccyjDmbG8NGWNSnbA+KrTg9IeS1E9ErUgjKT27nebzVQzyPndICn
HiwR4lhu5Lxe8H/3Piakpkhv15cuq8fmh3LXlFatFwyIYlFjyRywAAE0qGm2HbU4GGMfzA7Utf14
0ID/by3cepNm+6TY9N5x76WacXQ9gSoHQjzd/xMI/Nhtga1FW/56Ykedr/wwKEZZ8lc6r9Mk3LIr
E3PXvvQs8/gYDqDaiAp/bo1E5HE//JZVexH1EFKvLjNOUqtKv13bE6zKBGf3UyW2Xk28hkdRnM7b
YiJp4RiSA+DhhQdUg7Q7j8goGbW2N5c0wY/MjuOF1ZX+JKUvtcjy/tGqAYtCPWc/7Pc277qZNCv3
jj0lU8o89vDlBuIyywLTTBnxJmcAOqWq5J4EQtBTPvnna8+tmTjUfLRMlGUoJGg4RC4pzJZqQdgk
Y0ezranZwdVZpUSlZaDCurd02jOmPFtht+4vL7+rMJkNfAFIPdDE+W+OZI8ey4y4tEasNDB38RX2
mR+LqALaftq6bYYQxTipijy24j3588aKddtvMKc5wVHkddT6yxrC8tB9B0Q1jYFA6SMykyu+DWNL
vvE+vxvZyp7nJr4ZcQPxOE8JZgGO2RmXmjeFgMOGkwZmO3ONGQrBqP2ISbZqUaVXKXHsd2a0IjC4
1FNeOiuSgCBEuuDqnWkAcNZkKyAcD8gaxJxtin+UfhUnqmu4sucgEKYAqb6o1x7yXNFBZniyzZW0
6l9opVqA/RDYX6thBjpdxKPyUoi8uVZtoxEaXjV+lwDYDLGRO0rnfl5aaLl/3TdqUF++xeqHT9l0
C6rKnsxc3GeqZp9CZER3CwvD8/U3skI00bhSWSnqOfdZhDbaeqdi8/1BJ9ZqETIijiCe7uWBfNX2
11NjhcpiJOx5QIMs/ZjZqL2q/gCZOidzotoIwsEztwNkEoRBturD3luZHnPPp1hzoEpIwcYiaGcC
JkXII0314p0mdKKrJy1Cd8bP0WYKIMz06zwaRGHjWiZztYY0SkIZZrAWYjDbTyDU24ISXWzkNeCJ
SOv4acxJCGOreoUadGtMXYGePLwjNQgP47wC7y8koGZumAJ1HG1FHWm1KjPMBDaZ4pHPEGQHs9Rr
6F+/5vQSBQVufPgCrGvLbrBML9qS71IVfHQPvLQEJU7wCDMiGhHmG8m9qyqQ//vP1uvhjQv24QZS
HG6g3Y/QDVZFMSGsb0Vvy3tQIDEP/a6BW/NZDGIBx0LO0AibLWe06qM3o3FDuBJQjklVFwjRe9aR
I8C/tYzwLr95jzeXKmBGvURptKi7AwhdYgFMmEG61w5moUn4s+ds6SLluhIWm2O09E1zAmzz8w9M
zKUOE4izcnPZ4+Afy194HsHoS2Ac3I7bYTClZ4T02hImntBb3zZQ/h4ZJvo9/86vV4NmszKlmkc5
2D1KKGKeRYwr2ukhoUzyagMQ14aqW2o/AgHcwm2rmYysGJ/Inn6meLbZ548ZENUQDVMaMcDrkZDR
ByYJj4MKfz1BWV0ooOlo1ZiPkUd/9VDjCr1+ThrAWUEkzgadVz4zkLQJqfe64DGdHXFuFXaQAKNx
6gpbycZAAv8C2ipx+3eYe6qewe3NhA8VSuCcVeD3wmdA+9ESlrplcb4snvxi8FbI1bB+E11ckTkk
hDHjIOB/WOi1qInnmbHy18wKFK1sNYY/TamDoCed3eMKeRjmLv3aEXTqdq0C+y1F/fOFIV4yQaWj
rX543sRFFOFsWT+ZbFpwIlOcGaNMFr8qXjV9Xdn7lnjbEOsHvz60xy246KrvxSx09mSUIQ1kY0dG
4461c5ldZgeryDDYpEQQLgfwMkl0m1rtPiw4Srx1UkPP8XYG/h/Je83xCUrIOh9HW+2CIojpDFI5
24d2teD8nW7edQaoP+0FwzR3aLTYGj8aMGui3Ah30xY/omlzil53XOG+JRoqAb1GQiK9OAv3KMG8
C9/bITWv8j8Y1vU4M95exqcutZ3aSH7XJUir7/zpRJR0Zeoj17+wCq2sQWzj8RaufyZnEHfredO+
Xwxqr/grqd/vWQYIbuYCxkLRV0KovWLBtBHEF26873d4HI88pbW4i51gzmiMg76RS3GlUOYp0GjS
99Fk3RDEFz52MROPIaLewXCb8KQpgIX0pn/MqCLP7QiUDQ3rSlLR+g5gZdDueeoturKu7vsayF94
pWf34ytFVfeuaNA+zpwFT6U6yBytPfl0qQfG+O0n4DJA5CIaj4eZB9YzxSVbG5raDo4diQ+vCfZk
0wcmWgyZ53myApBMCGE4WbWxJo+kS8z1PaQ/EFw9A+0LKyv80S5ek4QDcCm0ejSb+8odtm8ty87Y
RnATLpijQqBz5sptUkIv8BDKZbi1aG6rpdWgTVQor5Uw2U3GarEJFNaZatCMYvJtOCERzPNoQmd4
SSSTgXG37vecLzW++g2Rp8gEkRnWjxBRUdv6zST7kA0Q9xVKSZF+cMBrnKdQP0scFAQzgGkGQD8Z
qrP6c8Ba5HgpVCNWI/6kxTv76S+dmIDxbpI4dvd860gih+OC1Z0Q9VrbXpd6MQ17+RBYFMVj/D3I
K5ifZ2r8/IHLyxVyHRDskjE7Nj53mqpFrum5E4GdRnkNY4h25boJBdAhK8dSpPaUa+v104jHTmv6
tDitIynoGq+TkEoCxdjcVobe9yVuJK75KA0/qP/BptHS6waCkUQg9VeM2iDxI2zpctlHWQH76Z0K
RfTI4v+VHB/n6zy915cAAi0+QiyJ+vyxztXD/ty9DPyguw1jKqHxP7UooZXtagIC18zfOjP9ASaA
Zd1SxlRpnI2Jwd7oyIA/sfrdGEPsedmJAG9JZuhnWN6eCS//hewZ0NvJzP3DZR43LmL3uBDHRpz4
rGwmxNHgG4f6HmA56JbZ9WUgaLGzbKwcBTgA9idGNvPqvHuvFZ1C1QvfTRDP1/b++flbSniepCqh
MBEPGRiepNUuGvk0m5hzng4OYfprcMu8JoNcBcS/f/Xzuujo50fOojCeyX2ZcOf8xU4Cn2zYQQ+o
uoRIWlnee+DUoodrtYakZUeEuhugUQTfWe0hcpfkgRBtFGvJp3z3nWXya2DgbBO9W5rZF8wcmLXD
cSARh2wXUAsXcuaKxyT6zk+Pg6/fAkjpNW4Kcl+LibW0Z7zeL2V5fqM1LRcU3M+o3vudsJ5IjRYI
DGxGky2ALoSHm6ZkrhUye8a9/Ve0XX7r1G4obGieVAAUJf+kIId7MVzGO+7qM0nZxVjIoOggHXdx
l+epkY+rz5iTLOcXrjrk1yF2vCzq2Ixgr4Tf2UVY0Lgb39ehlbGS0Q/DRm4lcRwt7m5a9nd647gx
aAs+QKwbTJiz1itJW5DNrxqojLlHWwxW7IuX6ESmPo6ELI9X2EdYHyc8pPwg1RznBJJXyNDcODdO
OPkZlD3Fz3BUoZNrdcMoknPpt/LxruQTSBtt/eTsOIv/ht4J8gGwo5+qdCsQ+gwj4mwazfnztVq+
7agJXRP9AEmZ2++QAa14bo1boK/s8UeAsRo6bSSbEILUr3Vq0zHiqTRNJF3cBf7htDgz9X8NLlY+
itYE/I7379+ldfAeh40VM/7jRsUh7SYWWUDButtSLRH2vGrpl8+uINWuNP4mWCYD/lA8JoISJ37K
wqN7OHsKcmxQ7GcqgsZ5wiKQeeY0KdHNf2LGpN2xdiqSSPIfgWC7uRDcagWXN/EyAbGUqDEkLGvl
qxHr3+onF1eZtjWoEzvoOTpJuMC+kf1/qGh2LuTnj/RD9V8hSlJLdKD4u04ofm/PH68XwaV1qoAE
g8JnZ0faqSkgoeKPhNiXQR0IFQQguC3AkcCVVG+xXWelZ7p1kj2kd5MC0W3uTaHWlhTbOldd9g/U
lThaEX8qiDhOv8ZIqqGqFkFNo8YyzREK6e/tRyT4tZ+mpLdl9CifdTtAFfhWneyMYYN4gc/kav7T
vET2Z0PF4YhxA8cN5D4iVDTrIo+PY4lchSdoZpq8Jar4yX/6ul0sfmGm9PKACJJDwoiOlU6m7NyL
vzgB1KFylP7qh6mQCZADXFUwDf3rtgfArqmO8jO6wC3WA37SPV2ALSymO/g8Ij/T41+Qi//7rv+c
QQ21AyEcVPTjKD9gyMAJMNJRJ44rTM8rZVyeOA3SkulGjZv7aqkzFB0jAreHXdUcSBHZYgh2ObbJ
U90X3rHkPZ2dSCiDOOZtrIM/vgnFIEd0EE9Uk34eS4U1oOXRFHov5dSg1LhthdWkXJR264IqWyTA
btY9hnIYGAnufFMSInb21S3wXmkTJdDj/ePFhFlU8YtunJU75Xm1DsSGCYfZOMLbKw9irCvA1+Nc
Ykpjj+eDPsDx8bztVQBEM+VbV56oJ1WXLqGesNUjgoOPHPKmUN8ad+/RgRxsCVcE6ou+WLvwEy2A
vAsGy5yZA9KOvvm9MUUD20r+/UT0AO475ybSKpn6wwA9Cp9AGw9jv/U/hgPtAV8pxjqHU1MDnxlY
pn/5KdAFdVFSatFnLp/mM0edvNXlDX1JXWw8fYg721PzY802QNWooA20Ct0C0HDYxyBk6j1UiwAI
Bs4CJ/VEpZzReThv0wpH5dFCozrT4UL4lZ/333+f+vRHkQRrPPNXCaP8jPm0c2kiN+9IEORSrcS2
VTqToJaUWX9GTzLNSfCVHj/ykMiHJRMSRwvIhmToeKbOsXaMMiqxDtOBIktTkdj8GJMnc66z4ByP
BlMUqfmf57IzqNI+YfGJSt7ubRezOlOtM55UXXyfK0f/3LMd67Ptt4wlpYd9EUtavDmKyxyku4tt
Wz5YfZfk4yp7L34QhT9a6/FSGOKLKY5XXPriXwhE+eJ5axqjQgn1oiZp514jvMS1PLEO8+XR7c19
DHrnxywyR8mSwB/nTEaZgMA3vx1JjGBSD2HLj9Wun0t2BQ+b6RxNWSv2YY62tiJXwahHPwbgdtLQ
zZhpXdPEw+ALq0c0PjSS+D8RmzGdwEi/NsxBvUbx1V1qcLWAH2uBmhwmMPMhouBX0+UHuAHKlW6T
tSnxE+srbxpV0qrSnJm9njTjuj3gGgwkHLGpSdIJVIIAms7dHrrNj7rk5L+EfukWmQ3PXESotGli
lMKjMsNX54PiT+AZabucdpjM9j+hm4r3SO3/n5hMYALVT2W2/uy+oO/vI/38NH4Mz0njpPX+N/y2
iz4ayrZ+3Uc8jfFgxhX9rgZ9kiHqBD5easijyzQLydyHbaxP68RAC5PPXhHMe+7WQW46KxS0vIT/
67P3cwwELiT8LEA6WKCmeVgEIB9A/AnFjqERekXsBf0AJuRVW+dO0XjybXdFCn+AzNiXyPCbgsx6
C9nxyv42pmJNjAVWpLu5JInqjZTSS7B3VvOtmDtjQPLwd5p+w+/V9l/DLtXOzBFvl3fqHZVIsJa8
xciC42YxECVEcqZKko9PXFyhWo8c/WkmijTjlkfk0PgWAZnUvJh4XsPHiUs36CSkALfj79gR4pbG
h0QUTNIwGFBwx+2JoxoAUrX8DBSo/G1xOSE+oLBKPpZ3wK5dtrANQaEV0G+12PdsG6gkPgz2f5ii
aji7dN/OT3EZQ+xG8gYDqKEKCokMeGhvUj8sUs9+GV7OK9IsmUziyaumyoeR8wXIn8P1vwUklRdg
G4mImJM3tpsjRtsTWV7/9Z5k6kRA8gRWaLrfbXWeKh0gL36GsIDwglf2NIzEja+Ikk1lbE4sHKiP
kqRv2+3nbCOzaVAvOclvUcrLrLvn0PPaw5Y3dck532Vq/rsNpKHCkUddexK8RJz3i5GKha//AoVU
YULblK8yo0SSp0OA/jyzFTHxHt3de6XD89DttDMs/5G72njE2YGrH5Wuq7lg+CubiWyhLzJK7WVY
D5lTz8Orfo7CrpOjqFkGUOaWD7JUwdC46PiXthYo9Dx+G4sC071uHqSL2A4vW4yjnpvtSVFv4D2Q
dEl7cZ5wyBAKWVKYW6pt6K4x9w0UZbxH+tk0BsldGrE+87szD/OnUpq8z9Pn/D9bNwb7Wx0IMMx1
Vt5hik6sWWpO0CPixeBTeH4epKgjZztr359mwBEfbcFbgPfJbH1YDT8dAWKaQBAzqX+edIVhqRRR
J2+WNveSNbkUkA7UbozB/jGl3hB8HbuArG3hzcTmpL0B1uzTYt3qfMppYrif7pVRkqjXTveoRkY2
/9IV8M7wZoqaDbrLpupPyrPnBeJqGcFuwfp2HyzAJjy/9qbN7wXcTjyhXQpi43jEqePVoO4zSDEc
6S2EQWDbDY/z9pxHhPHPbfwmoojBMgUsggPUHha+iUOI/vKHg4mFT6dBS4TIXlBH7kwh0ISgK9su
nnG0L+8+XQaAmtl7p1mNfzjSO9kKz6EkF2eIGYO4XW8t6yrX15Oiv8OWepCq5CVOXWhxpkwfAt7u
wnP9JPN8meYw39bcQe4Hs6snSQDb+2fuS6yBjB5qUJXa12LIDGQmyUx+09uJkG+J6WorvsgKtgS7
XFubZOX1IuAA9E9pyZlsVdzWiattcgj9UkYlIcWCwwrnvI2EAxL2hkf50nBxKgop3Qu5aw7Lg2Nd
Ctgen6gqRs62ud4qy9ypX701nfU6GcMrpPUUTB7omUHXImDdDs4Eoo+3Pc8R5cInWGXdt4KaTWna
fbsj/arHY2zx+SZb4KmWpYsMkQNjPg+5cxsjpz/Posm5Da1dtcHLguoPHGPyTeNnUfoR/JD8KzC8
AOkHbaKliVDthDnWrTX76iyswN846iOFNKF/a9hNzcU09kFh7fMNPSU7X1Os5pjVodi8XMkhzVhV
bC3WZfO5WRpzQTaG/JJ7JUq4IDUUMNui87DtrxlTN8QaacNX12OrfjDA/m+ZO3qEeOvco6RhE/fE
UXHR4OkSpHpXWcbKvVtPa7hxhbaBepFqagUd6eUPMAGAxIcUIs+D7v0jBwQxQEyA7ykaeQ9aPhXG
CidV9J8wzhtxdVduipcI1lGRpOqzCt5ErgqozqsiyBb/Hy3nQmCohRHtFNB6Ln47JeXSnm8Gkpex
ogJIBgu5xyodUgihiwfr5RMhAAMyv3uj3b94/4WrUlrlYuULGdw1JAN11/krkkUMS4AT5mar9Agi
TMiJcNd84NDvvJyrQjF7/c+FuWWXiMpza7DEBNMSlVz99Gs/wstDSX4zEZQtQzsNJll7fkYfvUoa
dGcVv+zlO0UQmmjBc1TQjL/KbnTdx6KovyZCiV/e8yk2kHls+7+fsrrAcRZrv6ErErlri44jucxw
7XSFu/eUBBl56nOMWHXKLdoVR4BMcDOEH1tsR7bea1ntW+iJy0xgPLDahxNJXF9xxvsUx8H0CpG3
iX9PETwiK3Z2srF9PSHAJsxdNVFs2JrfZiJjXvUj2mg9gEymzLbPcAv8d+571POlSRramKNoJKwt
RvQEf+ke5lrb4ErBitr0FwqzZNWTlN2iM4T6P/gVfjOwcNGsPnU3I87DslYMer1ZOKRot9+GqRHY
c/AmW3PAL82ccjwG+NWITeiaHpwWW8tommzR3paiGvGBuWGaQSrbzCL/xsYV4JImpM1h6rYQxyDB
DgmVY7NbOMNOIDjJWVL9PJK91PorwESVu3HyraMOFVHK5Ssa4O7qiER2u5EfDLSJHF3oevyx/ASu
Muk6O+RKMYHqy+6PiIfPs7PrvXeFKXKmdLqof5/0Ns6RijAC90zdSTFMHC8DZ5rzU3abaWYSsMcS
n3JVMSjJhtdUpzAD0rBuWqp0dK/2Pue4DqD/xdBv/Ft0Ne2C7MMOKvt/sk0Ri6oFKJjJy948IGbA
KTamZjC8wB2YV5p6Uqk68TDa9DbpauVO26+heRAUNNDP2qvU0ZWGxtbXa1g1qW8iSxahsspsTVrx
CPyLlym9X0Glp0lfyQj+VbVjZlV1gRmTjRUHazirgaSmsXoiOU3CrRaEy/gilyPpBdNoAaCjU71Z
Slr+1a7rp4e+UWsSYzFFLpp3vpZrLa7bRZPLyOKNtR9jjqVLzEGZa2rb1gS2MrLkCBxO6YypXfpn
21/2oG5zBTV4M3pg44B8qW3GGg20UNGOSRl3vegNmWg75x/VjANDy8xJqMpSms10nngdZPKcx3Bt
o1HWOjiD2/B0roB2hkXK/aOKQnuGqSn+TGM0oknkl9X67jMHUvT5DONr1iZS+kqFUOgOTT93iFEq
DWn79O2C9IJmLsQ08dNx7Sdt/6IC2npkBJrqfcDSE5oYz6dLrRt0y3kDYMumYXJgH6PziNtaWc+b
x33qhxxcIRjryFSJIrbuuBuQzeNPPQX8YaXH/8RhECLI3ZCr7PD4W+P8W7UhGvdGdYJytxpo5tc0
WZAQA9s/nha5Wu2k1p/J370Kj9P0KrF5Y1PUe3+zPLkJq4RIrE149c64Fpd2OCLQaPUfL65Bv+BQ
Rq9ZYnZY0q6ubFLW6PRKcUrBuy/uvSTu5ICVxTsbhwKFnm5+4Ywy7GUXELCavb0rpKgj2fr49zxw
20CVtdDtx7Uh6i1q1A0H5Di1ZAq8mwjT9SjRG/rbvSbtXAgTR8O46vH+R/SUq9niic3/xnmiyY+r
rFv5ZUuqGMxMVbMdKqbaTcPLWI1mSUUIbA6B/GkH69DWhFcyfWtdtvm8a39/HK6KMVVyoFWa+WN0
EHLR1mpDy6kk1Eh4OkUlV3m5cI7XsS8cw54f1uYffH0Uj2L+y8Sv4bejWnXjHohsvJRSY98SwJGY
tzvSQbnqYlKIneFlsX5gmgPnCKNu5loKYp9mOSIvFhScE8Dg0tUiihN11DdIwgzUZthaelGJfZah
dwygiUIb0nRnJpfUL0H5QWyzNbX9qZbKV6d032QGP/Pg0oz3YdXMk90g3a5+p/dQMnasj5OBRNQp
vhczU8PvD1U0zFFCDbdEu+JQSMUFx42wZxF4AcBAkTtZjyQrpWogLq5bJis1YaDG+UoNBuRDve5z
BBLtKdLpyCmhx8jl47zcofz/elT5grXD5cFmWHBXpeO3JaznU/VWe4YxtMmw3inewmLYd4NXv7N+
E6ZrgQsViEktVdkFGIg/D+lB+DF14K+haZS0X5QhRVc19kWy+wevVpEKrDVKpsZWHSHki7AWC8El
wCs6V9X9Q0K24pNsPaclikANoxHx0IdMcSHES4gOGTF8hM8tUV+eBodV7Esm9lHRTw6aX4H8b8Ys
uxl8nvWyrcvrvl3JvUGR0oKdhPyJMctEHeDc+auedsgXhtSQ3TnxG4Ea2FJ4Klm+NX5b+scvnDM2
4jsvyeemUKgT/wZ6eVHMST9GOp5I33yZuh6h39BmUaXf0FvlxprnxdC/LfDIAruYmcgAb1gURmGP
LLPphgaZt+XXGS6cDRtzMY+L5rb9hEl69szfRC1pNnfNPkTcw7NOfkud419yX85LKsxsVWA23+wa
IYIaHOVlFnH84fCjBix73L6qY+EEufqZcvviP3affYTXnavgzD/U0ILUp1YCJPe38TlED8509Uqi
YklJoOz6dLrTpShoHW/aKsuZ60sXEGwh/B3VuWyEFEvJZ3Ow2z5Mi+Vii1Bq4LOAN5xd5oHNn/bT
5yL8aNcTgoQsD4NL1bCHzZfsVom1ZRF33t5oRBSb3Bseb1Ww2ntDRp4PojVc7A5AzeYHUKEs7IKL
qkeATk6VDpFu08TxLK244bYxYg7upZQiYjnzGcFD5DxpSS9JGVQy6a0YojNjkTsevVhsZR2XDXn6
ylgvynVLdqLq6vuSX+VRj4L/hxccJtZTawU9oDcsMzsd0pi34XRUQKpgoJSmy/TYzkU9B52rLSpJ
vrnj+4K235V2T2b3o4tdqQdZU1qItKN6RuavJsNccLpw150JPGOHZ3JNPgGxATiA8EdMm8uWxg3S
LAxlBjdOvn6rfkovYwZLhK56h3ZlfUQEe9vNmeaKEMLmvyUBJ5hd72KnK2wz8H3iBy5BfloVM4Vp
xMtR8V4m4GQkNXTgme0wB07V+etYBRAsHuPBCeG5HGqHrrZGb/8uqtukkGvm7+Ve/Dfx9/cdVw2f
LqWEEbRADvfodl05XJZqUTUUbeLxAlHywf8aq8BY/ai11YxDerGvLmrlTcja+YpNjZUYJeYSICJ5
+M/pqmegbQwSjScQMCLf7oOMRMR3hoTYof4MP9HRyQOcolFBzw21FhnzYUDnKZJPxfWU5niqGZwb
8DSq8IoM0wlreesoPFS0mP1IXfqFJGX5S66RB8JgkpdhQppvzeD+W94xlJ7vQ68PuOwJORc0enI7
eQST9R/NiDVlTpP97yr4CyS9hrXXFPWXBePV3Byj4lzomb8EWvWzsyLN1xAo0bm2x5I581Zyyvkc
V9AzM5HJ3FzXwBY3yFIzlqVzveINODAjfxCACHFH8kXpZ2dTvjWbS+jf7HcpdIpt/FkL240gJKDm
nVhl+xR2Q6lOAGKNuvHmeHGD/H3YcpExkdFdySsRcjsOubupBtLGfvsCLLpCNfNUx3QC3uh4nNUE
36hfVtF1ZSLRFNAKGGpE4/XaboPKfiwpepIGBrY9YBR7UAT0zcfbdRAz379i6KIA2t91mpQ/rIlL
EPXSigZnbsh4ttZ257x10H9B9CyHVgXufnkTbvAtxk8XqkUIywyut3b7u2RVv/k6/iH766UtzjgZ
6G66c5Eo8HqZq7f1oWxQ246oOb2/lDgV48FUo9QEaZlFeYIvgbsJJqLNGxuSIQghI4v13jX5b1EF
dUzWskejv7biQ6FcxL3LJs9eBkqi5rcF39vkvrRxCmtFjfQ4H7HhKqKdWmtCQqYb4SPZZPK3+tzJ
VYFOEleUG7sdFzDHi0rcmN0uHAdZ/PQ+Pem7lJI6gp17zzVnvh8dzVviPdLNKFAnhdRJJdcmXxAd
0P85hdnRyr9vfu/uI2qGmfoUxREfmQG7jx7J5zFV+a8G5GwmAkyAlMrTL7zPk7kn+SiOFa/UlUnP
28BRX8TbvZnNXpaoGwRh1BlDRlJwNY3dt5fdp8MnNYMEPAnbxkc0Xe5BGAS7c8xnbFiDAyRgiIei
NgiuGxWLQh5KCeBCnnhitMsTkPf7tm2ni4W/fWz60Y6ucf/NcD0tzJdU/ukiJVH8t6yMdyVuugaJ
ux1hQygoQl66EzdnORsnxg3UfznbAHCTIhH3JW+uUdYsvSBntLDBh/KaGhwsxDTP5ncWvNfDg7zN
BmDn7aSEdZDKYQkA2Ok/1qvDWWoT63K9aqBs9eBLMLD8id4DEAmWYoIXr1cN2eKNlP8cfXxqF5q+
Zx6e7PjYmomZTGIP2T/JtvhkobjuVpzXlu3I+aGl5V9JCKv8SQ+NJ6+Fat4/47cg0WeTeW98jiac
lwgo/nxu+Cdrl4vftBDu2skCRUOw16N/o4I1KJTbWYX2s1abOttRu2tpW/vX5jdt7IfFE9xbWAHm
ugR00ixCgPxmfvEKclTqIl1gZr6r/pnfK2zOJGWIKiznF7cUjfAI298CZRQs2sBHpPxgglCzpAy9
QEZR3MWXdefxzlDhXCOupIWd1PVkMy4YLgIJoLpPMmMnbjCuMsAW5AHIvDjYZSQopRIBSxiOQxv/
iIo0xd/j/aCb+Wfizy29U0A/x21Zc4xdlBDDqxbOjoZNmBAEELQns5/RgL+BJQJz9i9C61xyIoij
3bKHxV/rVK8qyXLID+3fEwPk4fvRBuRJyfGSjLs8gMpx6wo5VOsK7CyyHoUhOo3AX5tZeuz0V2Vk
L67Hu347ND7lXyicIazI44iyuLmutqt7JJ/1DreATXLCrxezZE/aHlNNu+A2sf6pZyOWPGHSC2OB
CsgMXX75W9MCs2kGsnZ4U6JlXCgE/sMm99YYCLDUSJVNOmfc0i5geINy9HhSQ65Uwu7JQoYfp18b
fRNCl6HaIJ2Myi1/k3A7viwDM4Yq03Pt83Xbk3vNhKWO11XV1hDGqAYjQy/5S2Pj4+6l8VtV9owf
NnalcfFcHkI1RLClx8lIrfRdnjtw1tNr0w0WbjORs3qftBStTyr7nYzxqpkTRe5kL8X35bDkd34P
M2PfOWE4e1K8b86OMyrnXv+ah94pQk8xf5SzM9mwdQDqxPiyqiRM78LhdVQxEpHM/Pem1GumM5dw
eoCeuibcUfdBioUM/bWHaN6fl4QpmwysS+risq/wy0viltuW0+0ALZY/G+4PzQQw0s/k8Vc3HVBA
DUPwIs0rBpmY82P2oejy1pjj+I9DYWAmUwXZp4v90lKRhA2/bwTQ6vADDSo5NmohnX8ZW3D2ydha
2SQ5AnAAChW9B/oCbUci+KQOhvZgeDSNJITrlg3XM2x8C/5DHnUKe4qkdrrKadjewbN3p1UsbxtQ
z6s1Z4sZ+i+gyTOlBn5TvZztwe+2jWfLDgFk/4R3+Drn2ugQI8Xgsng5hV2fRTvetWhtB30xOwMO
JPHt0A3dhWnMFIjINUHkCoIe43L+K/P9IP9H7YxnXv3LihDhD3XR/XoyDBxqH5J3GilMW1fualZ/
9X/EN3yvuoFirMAgwGeGOEXToqi2DjgNtCnD9cOrNGdKGQbw+Pv2CLw14XNE7tP+dqxFRxixyaPx
35qUcRtlPqnlXOxWO2MO4DhlhKC0EN5ClLselaIYu+1IJxMkERsuRUoV8ske0lv4mtoqvfh9ak20
g0MW+CCov7udtck6o3u1F1iyiXp1VIHdODMMSGJH+wOvUZVSbGko8UooaLbj9JGSfag8JNDqGVAl
raGJR/80WLfJ6sRk61rAGppxqeWci+HB5Vr12ZASLtxHBu2B326u/B+tbClUwcLWl8bhQ042Tg7i
TXHoHHiSvsYvuIuMlaWID4OkkZg3hwRbOQDAlHJWOnGv2rt7c9rjEHAnDYKxLgltI4CabuRSHNpl
ReonhOBh7rz3RaO1ZIyeo6tcAGS6kmTNiDEt8iACgFoEwPKiryZ6JvIY4/QdMYnzeE0eOMpCnOuq
Qw5624xvYlQ+xFvkBi6QQAZ8RBwF+kANByhl5cZ076Bh2DnqTRt2DWluxdSmV+tJ+Fk9o/q4Ye39
bmxG5gLcMEPAzLfSIE4CmSCxrHtyG9IfKS3GGcdFj2WaOQcbVDaS7eJPL1MxPevyFqspiNmOMSuC
07XHIHpKSAhwvsKykMmP/Qit+sAiCEg2QpkGgPKZVj1lY75JRqXQNyLgxL2vmBXznrdy4mVzEkJJ
GIpD8XqqwG8vtYQueqncE90IMIE59oDXaktjEtOOFfoSYQIjsnCCpSU7jku+LkResWoKv0v6NhQY
kyP6ojQkwWkQ9l3EJClSeRJd140wloEmmN/PMPPB3Te7ugAAtojom5UtXvmNgr64llZ/2jz7JUpd
xqw0VhrKFQmMV0bPt2sj4+HuCVpWNY8qzORjCCRF/3mFCZNlxTU82lbng+yO2pKTSgTu6peDJhOB
7SGKww0o+Zl8yAT+gez5u3y00sn618QcNLrKVVNj7qyG0rxSOFUR0PRZX5nZI+9IxV/B3hnVQJrC
ujV7L/OVbHwoTWFIxEG0tnC/N1d73X4DOqLqqVl4kMIo00VmQuXavXsFMTbqINNlsTfaKe2ZG6JO
aqcjvMeZwVsBcNBt8l45R9EvJ+1J9Q43hAZX8c1W8MwKf+w51LeGZym9+9cJn1CFKSJCrmqfz7Yo
WL86PnfLeV5Zl95YuPejhsMjcnfKpEzNd3hqrGQhEQwPdl+ol55GFNsl3PkKIA5+YyR+bYfccElK
vtslqpwrO1kcxfz/K7f088ppREdQYDREv0oT9+aFgSjuhLID2hFAr01luAS4rX8pF6j/g9ydiI6M
7HnrFzAn2OpxFz3ti2/jRkoILzOIVtjSD2VNB539sveCY+1i6ohAeDHMrWaiPgHtFt8FDVcZIMIE
aMLtkXbMJssYNfYA8N3my7sRG3Lq9E0VxLE6QwChwKlv63f/wskkXlTAFMD7zsrT53Wdz4Lr39lO
yS7EZ57T26tk/J0v5s3D2KVLd/g2N9N2TDVARYsPD/P6Bd/pKZbRw3lXX0Qeo9qP9btpbGKtg/tS
+IDkjB9doNbzAy8OmPTetQ9tbRK7ab+HhSKL7TmhpaHDTuoI7ksPkkNaQ7TbpKGfx7LJDpWFQLgT
J0hXZg3FWX5a7xcTNn+OBGANl8juAK+HG7kMTMox61Ib4oZXowjex1Oze8L1QioV2eElomsurI1n
bguru9v7fJ29xtfOiajzTpE7FH2QJITGTpU5FAOIhvFERmyXyzCJE+xh5CSPco5fYFfFkOsofDB/
sOmr1VY++mN7LtkiqJqhafn+xEsQoxNE3PucKCes8WFLDJ+s4eFo5GDdtKrDwBrFWFdzLsXP8OEd
+uM56JqjQYVijY37daUebAN4DetyieqgrmpdRLnapS+pTQPGwqjaB5ugGDEbtSl22Q2y/WKmru09
e9Wtf+qisupImhF5hPQxA+EnItMAdhTIZCP1sxnpZDxKgDlU6VIQFjnAvOd9vcMNaJ7WfJ/albqS
M0Ejff30wE1IkbLbGMYehjdvDhXHXL/MEuCAubVonaUUk/YjZVyGPkSOeKMeHLZKomaGgS/xqK51
aH1VR9em7cvfY/17Gp7GvcNVY+tEHFdMAWfMJaw71g9ZZXvkT7i/f+WyOH7jyRa4EGXnZ1+GFPae
Oz/bsxrWqYVUnxbyp+gUvCYkU95xSkYp9cJ2hxum0AJDGE1RcV6nf4lyU+kAFbtcLgfuoetJux6z
SZzEffVFmToubRPiyyUHgEpIv6E8v2Ec9J6aKbImAOnKPHNFi6AbBRHImX0kUkFEJaKf8c5/PEfH
m7X0DEiMmLRfpSjPqYiz++s+fpP1b13cUdoVAg/TEOmGr5wi5h2vRUOtt/eg2efq/Pj/pahVTlu1
8rBekN+pjjTQXG84wmLkKTCXvK0CX7IsVOZ/mhaDvzSdsAd6jeSzaaOqHyazjDcc7FVy8HhknjBS
vWJctzoZO1DKfi4X4YQYjRzKDVM/y5ilad328cXtpFUENLuNziMZmu4+dKWLC8iK/7/7ebhxeVOK
HlqnlTHfllPyhJOX4icLkE+StruBDNvTOcA8ca1nqgHGws1theUyOOeHKCDtKUj6HODwYs2maxml
hPBunVkmE2TbCMtC7/E3TM8enHNDcbND9GkpteK7Xr6J21y6COnPCDqPNNntaaOd8g1FhcYz6xKB
3chTypx04CWerOjOnPGxJWteAesy5IPL7w6lmPP8kMLgckiHkMalm3pGtoV1vWHi2je9oEgbA7qk
UMx0Zv5HRWmCHJqy8U1RSXzqQm+6Ce7LIn8qGqymKdjSdbAYkLy00vD9mS+j4PWxiNnPf1XFIrBs
Lsbmo5x+RBGc5o/FjfEB0uFxBFFTVFj0yBIBAI+WLR6p3DSrEYBBskwBYtiPG+ak+rXhLPLp/Cif
TusZ0t160JiVhVSEioPJ9h+NZSvmpkdcECVG4rmc85ZHxt7NBGcrRfOi64cC50zxzjLH8BOodq+G
Na2/L3p1UzoNKtK9X+zGtXk1uhWO6YcE35tXqWsBkVOy7qPLX1an1YHCJkao1zOao763pw1jjLOD
edm12kTveeZCdyEi65QArKbxcxw6FePLnxb4UB6HmWPO5Zntda5aWu9nCA1oxaSA/v/8r/0h3KqH
eu+1YHb5wiJbl6YYN6zGlrpZcnAK034er7Yyz30/as2FLJDH38K/VLMMHK798clifAyJluWFEkLG
KZv6e//HCll17haD4tamIWJYom6MelhqU4Xsq4HMIcmhjcwKhsyvZWYKlZvAjlLaJwqzC9i/Dt5s
9inBGjf+87nPHh2MY40eYpvyga1dNnQCxV0AB4fQq3lVkPddLKL4Ymwpo/ROuuS3NNUcehPMngis
7GnWifS68AGc5BnwCnzZTAPGpIYEakyHiGME4YqgXuuV4xwDpzDDqJvSOCyWdQrL+BPUheSb1Kq7
WLf5lCTAjrbeOYpTyFvxS+8JVVt5IPANhvSlteo4LdGhab/MlD8DKI2AjQXyEPZTjeOyK4fyQopn
erxNMGPP0FDobIDU8NSOqd+zMgmC5g71tuHg8cCooHnCfK6M6kKMRg6o4HMejJ9YsxaWMAhwQ0iZ
J9S6EBWcC7IotTSzeFo9Xp2xyxGL/DuEA3x6K9zjrdGdtAkyuQdHxs+5MYjsQdlaWGRM7PB5Ekjs
yO8T7DkFYeXq6/PHu0xyaHqJUToP/dIcrwo20RwglJPZ0GzassDoFb3zyAiPXOV6bSeAaqQe58jS
my99ljBZIeo7VJXNtiXNmfuhYXgaUfUbRZyqJLEQnNqFrL1bqc5XtkVQ79bqwLUYP4t47b2edtvb
ExMPOpavf5zMNKjscHMmfebJl58haw/numxtSZtXSKpoqkPGBcb4N5lJISDCqqMgfsREPJ/ezVzf
wuyON3XuL4+PzL1u0nVW7vSC41reKLRKWoxPXoigmAa4/bVpOYiuQlOtvOOfM26OghmxelcpOWB3
g8L0BqVFFRU85hOSeia2KfYzu/MpoLx8Y+9JxaRT82pQU5+Mf6T0IjXGFN0yTVFwmoi94BdUcyOW
VA+vaPgubHWnjSEzgnEdTZBeSrJM9cp2ItyaKPeme7mGSMNc5DB4GbTryf89SuOlwzwzg2Falwmo
WVSHvHKOcCnZ0w7G9p5HcL6bNXJtLoSoQM9gBjWaYEEMYcxVENE3Eo46FNXrC6oyppEMQ7ByJ0Rf
BFJtaAodiQBVp7LQuOzSSDBc1Fbq2d9sfYEbE9faKLh3TtgUrTKE1mM+eNVKoQj74QPAUmku3eXa
uk56c7PNOG2Hvhm+F1O677qtGycBmlNKX2Cge1c+w5r3bS7TOgPz4V7J6xEYF0mYlDJ8SjZLG3h5
I5/Qv5KBONFusuy+1lpVP+H4LRnNd2/vslSmnkZbgGwKLtwqqQfYVg/lxyoPQkS2KFkstfR67uqN
qwIsQm/rYMcJwwGl0O1QdAVkth8B3QitSEe89lya+xRr8N42YTqopIsV8Uk2Gv0z2lwkC5adqGOH
+tKRDPFL5+2sUjq0tofRxWRWAvvyMsfQqs/jwFLROaaegn0sTPWqCoodqvpRh3uMzwazNhxMtrRw
Fan6lL85jfCCQG6u8GjGwWrRaNxtpgSihVUDtRxFAscfYOOZg3fJ/JVNGxmHbnolUhg1MHtMOW2p
QBTMD0P++/zhlqyDEoTCnRAjKpRP3nkI2ZKRxOybdozIM99MLpsH0yUy3hRkzzUCvBcFGTEx11CF
q2MBe8DW7SV/PLJs5hQZTe7FtDr1aa/2b+iZba4h9jjQSyUCACIKq2bzzn2YMtoukbe0AcNMURDv
1C2JO2MZOl9H8tCREWpQtlSBdJdCxkNya3+lbCiZl8l5/3BbE6xeCTE4kIivX1+IT3Hcp0me+OGe
GO3KAtMiMBYG9Olb81CMzh1zMB6VDZL8A3PZ8XxODclCmTFrYG5wD5AY2Nre9o2VBbvri2J3s9dy
WVFnc2XPWyp0teWlVPFweFRCcD0T9CyfBIG3jrAOD+Q1rF5kUp/7gaH1z+V2sw5iIatCCiJxxCxv
3/K+k3ibv+dbn2pfOYGMVTRHja5N5q1T1MikktupqRum/bQEmVBHD3C6GPwVZi4RHqA42TEvIjiS
bD1iXBovrouFtkEKPdj5Onu04MrNMQytqS/dptF89XNUXMlZjLz+7LO8AaVg5OuACY6oLzE9R/zP
WI0jzrT3iZXQe4NgseSYF6/94QzYbuh+cAYPNd7bg8StoWbwqe7z27+4xxXHgNFIP7iewSqF1ier
rEqbkWPEZrX+aYMbpDtSodb1LjJhcIH9v4ThEWxwxNq4f7YaAQO4qKdGGD54f37KY3rifzyEu+VQ
RXyTAZt8JdQJ1vi61727fhoxaugZCvu0FBltnrXl+uotbu+tcW1VVeVQqsILccf4ysgZN25wvxuE
Qh1j1vCimpuUEZq+D57CI6hbGHDp08YUHjfIjkzyp715N3ivQtbMzgJIWxqGjLy+dIafGs5yiXZH
T1+7g5hJ6jBoeIf5TruaQIVva9qoP+qLoWAbz76Zi31BAd60TdYM1Orf8hm4RLl86p6NSWNzxH6M
sKXNRJsJhlz9fS4Lod4Wu/n7PGEVC0Cfgz4COOFppCwChQeeJrIoliXalL6ahXbL3k2cIzu9LKTz
BeljTbxdJIFQJOyelTtyxEhqsVuz8zGMxvAOaKFng3RLL0e4YirGz3yuf8bTNQc9UZUDHd74MZNJ
arzSfQpKpyJ6ArAEo5J3vVaw0rpq8Lnq3GNVYcxk8ohX1vt5HKQTy1vn7JrI884Kyz3/wwXr8yhF
i9MQNHjggwenHiwDivDtJDiQ8WStc7aCFPjMjw/dZPzwWeHubdmMmKz55PTrQ8rvY5p5oI5EcqPA
oFVvHVHGRgWK7DAWyaV/PhfzfFU95g5sy5jjkIPn2JWtqniqrj9gBD4jTJJfqfa5wtzXs9SyoJcr
3xPSoDq5yTnIsYnHPDUwT+llJumxYM5YzeEmajr5U55qgB15XyUxXFfLz16dpVF/cnbiz7cXTFub
kTHe5O+1zxLqCW3lFM3EBtrhoNfk58r7MJTNg9JO0mKkKQb6weT3WBRPyZQHj/jxsFCxo+rP0QaW
CEUxXZULZ6Pa772RH/0WzvMCi5EPohX2T3TyB1/Wb0WeAK6PLY56h8doLCsfWDkSc6cf70/QnTsQ
QP3Q11u6lx3P3mfFC45HYNJXEduE/N67geairxD66i7+AR4X2YnNm+I5Y7NEJHAHZVBNZaZ/h/qJ
Q18pFrrEe0jFJFs37IfCGN6K+iFqrxpyf6kNVm74Qxsi3Ez33r+x8b68BeJGipw6I844DFurTqmP
u61cSdmNd/CScypCjp4W3a55hxAO2czNvLIutEUhbqOL0Er2X8gBw3asVirzDP4mN/NIk4cE5yt/
JVaXYOrMP4u29pENkn7nPTd+VrtMOt3sudKTcyBJF6G9vJfMcfofzX/DAYnfKRrnVluKmHPKhTT7
eC/MP18tbQxIZjw88kGUGjteCu7t/XAJitml9L32SCNpPFBwInBoo1VWF9q9SJlNrcAsnA0bN9pd
c1Ra/QfKA7rqJlKsHLGAEmyH+7xI/NzRc+JHBcXeYg9Nw2AFaqa9c4JNq1gWoXRQzj4tfZD2iwQV
LTsrLr+yec6zYoOC68A2f1/HpWptJqKeEho1iAa+fatXEurYY0SIfvNNgZ1XxINPhyg/MNFToj5C
VUPbYS46SmPMw397jlbo0suqkeW8awpveOA6Ohgu+CvLgMrzq01dAJp7C3fjvIGQKm0auqW523K3
oHrHLkyHNxoFaAxlZWxAC0gBY3oxXUTfuxHDxiSQ4mjrOYXPHMz2fN3bnWbeDk+v/RG1CKqEM+2W
cZB8SGLiS7hvlA1vo6a4Zos4BGIgrjAK1fYF1K7XnVqPG8hgQmg2Rk8dV3x0Hig5gfz1K3FWOMX2
D+IBt1FTrPP9jfzIEHNlyrBAoq+ReSLmE7WxSGTJTy+W4VMf/n8Wh/LV+ZVOHkIMgMM6kR/+ROKx
1Z1JegXbThvsBgcdO+5YRWpIHVR5SEELngvF4Oz7f3M1cew1i9aXUv45zkxFjO2BMOfeMnvalSzu
XI7bbVl002/RdxeJ0LN1H4b/i2ER7/NM+sqLrcRyBMx0okZhnwIVLr3hSkCPRDxPagJMBX8pqQ/A
Q9vlxtaxQnf/RMrobPRoKvSOKXvmA/5uL+eddQyCA1ZXctH2NrsnhYY5uqJGAW3UN8xy+a6rWWty
+GBXcnn2lgSj+t/Rgc/VaP4K5QQX6Pwld4b4ZTRApVPoLv/Y/YFHmTrgi31PDhXLAgpKleOvFTV9
FEqr1w/g4IxfXjWBoN6QdWfIx9mpq4yrQu28FxO4dCdczGOZ+H3k7iCmMzF1NXGM1168TAyuFvOl
o8ezizy5/ANi152XHzI2kUa1MAgBadFI0+NuttqEmXgT5xqOT0Gq4pQCh8HYUWK+ylRIz5FOoaII
plXA4TkrlRU1FELw7QoT+/N52cAZQTI3qch8gvbugJx25JLyt/1U1c1JCTUp+3YlTelRtYunPGcx
rTyUcrimK0lrrs/wXDIjF75oY/bSwPp6wD9p1NhQkmzzJglxjk1drqsilGzSYiUMnkLVo46ZWKzh
1yzbZOxM+fCM1cxygXVh0um+L7ARTigFd00MEmSwU3l4pGasLcnkVIrz0GnRmmhVg8RiWM/W13f1
WaF3plJ7cNLKXFc4q1Y1OGwq/CB/wqrPM4tGJBol3/fcwyLPNYPlNSZxC+X+pOJLLuFCpIzuVeb2
m4H06LSi+M1X40KYIrxekTDsctW9SixcPFjUhRjFctxZ2pZbc2NHlyL7i3ZKZVGqzPCG7R4LaOjI
EgVcHTaIqYMzdiiG4iC/DA829UkKALbCxhxos2oepLlqWSu9dIDR8SHybzKD4cp1WJL1q/FWA46x
jKFcYjpLX13Qodmqcrl91NPjpftStqw967Bvm0bQKzIIvlFSEnHU3ZXc+y2qIaU0jIess7ufTf7J
dnkbLbA3WL2O+qu52ZJG1aJCdV4WawzVkoSqaeS9we2vtD+5JNKuw6de5sQZT0WOXowuWwaselpm
P+DJJEGhjcDXSXA7w7DMWFdo6Zyea6iGpSGNogTTECnUSTP+2Sj6evdAbIVk46T8ke3J8N+tsUX7
OkOTvY+m3XZlPG4S5ihs+Kl7iJx2Im3II6o2QVBmtPS+rhOPQAQYLTIYdNsz1upkxdUNBW92kQ5L
PJiGZMnNp967RECHRftu1oiopRQpzl/+A0BKXXz22bub6W9/atbq5mGMF6TuiJS/fWJlbuX9NlsZ
dzLdLJXAKUYNXWMp3+1UinZsZljCybqBpQQhFPPwd8d9eJRfyPWqKozogWFRWqLcFnSyHE47cHLQ
Y3gJpWXWfBNkuICL0AKaE4rSB/u9pWy0F7UfmU72PU/FITOPtQ9XAr8w/nZk8iyd/lEiqJGKnbwq
oitYbClTU9ntxptMAczqxiUTXbqFQIkj/OsNF/1NXmJOJneufslGBNUL6Ph8bI/JmdxtDxALbzGu
pH/jkv9ugJUk0LNsiJC0E9jBD0szIjv28mGkCwbpvRN+Ez+o5gfGa8huUZCwdy25fExqMZNY3cCs
gYKXo4+La+AqQR7achpFd0Qr6XwVhNLys7VmTuGtdu8FVKE9r0GgJPdmqvODHyuI3+zB5I8ojevF
1NvJ4M6jKbQyoNPv7qhGbeCV16NXH1FtcPPFz4DZTOdVD035jHIuafh4xtI1yWI2nhT40P0m99Oh
Ljwzy1VY32f8zXDGdJKjsxQ9pd7IB9WcqU4+noviV/h6mx9ylkNdrkzRa3qCU/XrxZEF4quYlVdC
h+HydsF/OwYn5XQffcpPcyCKeTb/k4EfIlOv6lkJ6f9JTZI3lymXTincbIlqft9ppnidga/njYbJ
aZZ5MbTfUyKWEY/DDkli4zNgMUpdpGuW3jIL8pprurbZG2O7Mjly53ecf45TH6W9X5ZEWXJGVvD5
ByMZXo1xx8FcZ6qXmryg1dokPodAXJEXj1+HDl0jBXRO01cBehoRhZVd0VeFmArTjcz/cj+8nQtJ
nb1fIo2MhxfsuNdE0yZXrGsUjEOdVFULHY1zaQrRrvwUrh4JfekQ8YKAOCzd+Qj+0yf0H81I64hZ
ZA6uZvn+30avsPFWAiP5j6SQLse8TJYWxy8vbUviaQNHKhajV58ax+K4fqqWYe0s+WmWSXMqHJ5d
HPFfzZMeCaMqVHLa69IUvaQlWAvSmm/AhgKWbhIq8z0a7TW9iFIwZ+f+yoD/0XEqL+1ib4MhLNsB
XYT3N5JI+OMkIPv1quXhodNlf6QjrOlDgjV0j0AmqR+r+il/aC7s+CZCHyWTNykPhMgcrH5Xv8zP
YfOu9v6DROfRscyMRbId2vfmqiTxN3SNm4H0T+NZKLnDfUAocyLaKppIIFu6OwhCpylPkJ+MKzjN
61bRTqNu4foiDUUk5fFk8QkherqKQN2ebf6hu5q8bqdHh6q8VZX0bRDLJfRfAIMRKc3H5pGhWTiV
slyr8O6Jd1AntcdmGlf0KzwLzAOwFoRqg9Kcx2uTwvkIHEBxbToCuWlbQ/ly/wPXiujEZOrPx5Y0
1yu48pUyFN3lz8rAxgczK0gRTlJ4lD0XYLQHcpLME95kEjWljuhggqkhDvSZCRSo3zmtUQ8HjQAu
6+lSLnD+EHNzW+WinlCbve2oZTK6ham5khkVj2ubEQObyOPHzbTRXqT6N7VS0C1ucw0nlsO/8gLX
1K/Te5FfoO71t4XrL9n6LlLeKwCWt9zL9N32mcoTq6IiNoGd8YE83qK3FOcMYIFcnXiH6fEuyW5c
oUVUs4cCKaxNybMkoASs9FoloovgCXQrDKZpkmOXzQcL4UAx/YgAvkXfWbz/mH/KUz+pQTDfC9Wf
qPzQXBRHa3AOM4qEML5EH7LwTKAOExCFtKyf9ITQ+vpMsZr9xVsIYwiori5ONmS0nnl3nOanBG37
O+P5H0MyHDdW25xwojM8e8Cm2Omw1r/FOdVM01UsKwJ0Y+k1sY2dWgwb2tMeLUSftIIu5D2cyVo+
eWXyECftCUtFTt4d3lsnnm7S5Lzh3uDMTasUWWuurmbVsT32osMFn2ZY4JwtrgI46XKnxK0euWXY
NBrguTEy1Qsh6MVXCcwG4RLpVyQ6xg4xh44w1AVgmSsgK9bBjK0DgOQPgqrb7o0iOQAO/bXS1lDB
9Q/TwGWEEGweFCvlwhAEV4NXoCCTsoHK3VLYuFCFr2LBM9KZmIy/yiR8PNo9zoupEy7VCFN/lBBa
8nFEvrVR4dxj7InZYGHGaBsm3LhKZWUQFuJG3vkXYrjL1Ofr3o4RePqKolQjWink30+65pmCcG5X
DxtxcRB5jK5AnuqACE8RGl44UJvzU4g+eMolobDK8QNU1S6Kram3tjpVljIzDuT1lJ9ijKQg7XVO
Mfh6Q0B7AFtOu6e/VcchxV2lfEloNZDRht/2K54wDrXtZr9j/KoEDOMIVedAA7X9hDhi9ep8mV6P
JQ8OauJie8S0ca0tkwUoMZ3IwK+Tr5aSKSKqRGF6WqGsXEaKYk64IBK7FRGRH1/V/MEcOM/7uSuO
1mr+X+nzs1TMjLDTs8Hho97KWQgmQF2XdD5ZWEOhTGvR0yQE+fH0CODBfpBU9FuLrzdkAGMP/cX6
F+S6wIZseu9XA76qC/kDkMVMInppAn3HLk5tTPxypJ1HmVB5pjD0i7m3ucjKnDqTJa04lgYeU5k/
IW9eMg6XWizEYV7fPTZloYq79BsgZftE8iEiRjs7HoHg8fIrtoLt++jUy1oOUxdLyWHd+BnYG2wI
x5CxUf9e8u7WLCaH2b8B4rYjGBYxViiZvuUf5PyBbMbpbOvvRwKrFI/wgk1t2osFUoN5LJWKkmtn
ZMV04EFRJoDcTrbrpWCHhEHrwDGzeW0z7Y/DmYLZ/4DOajWY8KMqF1A87LvI86edfAIe2pis7odW
BLQTVbT4LNlV6394zDopUe3eqWdlYkHWsheVlpt4G8YQQuIVlacTi+xe9XBflVm6GW0toXA6ghz2
adZ2OSr4ZlA9W7EFCcS7AlL6412bYtz7Nfh2Qrmq0YOdBtDJcUtukqztMou5ysOH6yiA4WfzTYyc
TGsrvtzREb9UVEfLG413HKOUnAIWCQ3Hqizfq6R8Jou8B+TRaCSHlAiHEDXAc3an0Ou+R/jK2Y5z
xpLk5JJ7/xfjJzHqAqnyeDliTrdEEaafh28IujxnK8802XBa9mZy6buOKHJqmS8lRGfVwTgCzd6N
Aj2lZzL8zeyC07NoEMfKHRc0dgVgJwmkpkLYb4ru/zlBU/QNiPmJwPURE0MEgTbwGRO6G/Idzutm
UuLvIzau/ds6DQ3KFmD5RNDDLsyUL09dEUN+9FL/T6BrlqV9Dko6GNZmweQ8mCZrvcF3yArM+D1u
qL3eJeZ49PcFMhmZ1CUSPPjl6Ck/igdccWSe9pG+dCU8y9+gohg/JEKXpjVsOYZSxikGlQFZ9V6J
j+6OdIGOb9siRZa313GpZyzsHJz/CNpSta8OPO213GtUN0ll6I+pfv6UTRVVNaivTLZ0Xin9sbRA
bzt8H2zJ2qprbgOl79WhycXCIwgu+f2cCnPcGaq/OXy5a67wA2nAl5n3rwyjtUQLa+quaGIezVqR
WbP09O6oy6ORbsScH/ZfQMPAybumaypY13UZPEqCr8hTaQRhE79hzEzgt+Bo6S12bfnB1S6BsL6m
T11MsiuYCHopwZyyJqg9ffDXU/eRW2BEbQvMn4wvOi2haBVpk/yWWLNDRkAXQicKG6z98+wr7mZV
jdg4wSxfFBUScmDY+eQraTGUKDH9/QIDFMjUBFDgJO4IuRO+6OpmGA1QMwPhFGsz7GcwD/mAPd9t
Um9ke+e1zf3uAfsMpB8s1LKYOn7DIK+O/o5ViBBB2FkT5Vb+HaxdwV3pyi7ij7/GD0eGLiCh9P/C
H+Esfc8yhbwIZV2Xeh0voT746ejnGSPjYXTSpGHGH/9+liEJq9dWp8trfRVxlUfskj2zsHRLpMuv
k4bfXGS1GfUZHVCvv/kh476kcsrn8WwTQZVunrlMLtFOyxDK7GoGs4UpQUcxX4CP3EU3CdEoLddl
y1R9HE6rAdHKIsVP+0YMTkgc72Med5+brSawQ3jOevz/UUtfViPLO4eprH8cvZIo8h2kqy8M9nmr
ABSk5/sb+2348V92UE+nelp51Bs6sCwdje0CFMd+QowvCG3kSsqL7QhQUykz4qVjaiclK++PkTOi
i776wvZZPhmLmZYBI/Nxe7tut+GHC2bZT3Pt6b7GmJ8UfyCYV58CkqEiwdBMAvU7fYZPMmzdhZGe
hH1DFAfdWY1ts08gDx+TsfUMRmNQko+isPQ1XiSgD8Ycf0Ow1ZgKwevUIKmzd2uSGKSdmNM3MyZu
zsSLWoSHcqI64Ah0JWDS3yEELOIH1D6M2oUv5H0/qxeZchaJXrrReRIbBtpT+Jv5cB9XXNlKkXSI
GnKONMUN94qLfSkZYHsKfNkChd9IEpAK/ARbeVkq1pfMabkC7aQaXb8zutzr/LcfpUFI+rb72cHG
xGSTgfVFkDJTtTd9Pz8oR8ldaL14uey0pR/D8rxtHWXbm7V3cIuxpefmpdNSxsk8H89Epf1agrgp
lOQuyh5PfMZesSjrCIDwRjX0v/u5vZin5AoOyNnUXtTXS4ZPheyS5GmXCmuTTyzjROwCqwEfH8uV
NvptzuJv53eUJP0q1O+GsuCpztbWKdez3gL9iG7X/1f6jduuqTmqfBYXrk2fZBX6xF8iGnNFsekL
9lqQqD3hD2kiyG3gQwGxAbNmnuE1zQdMI0kgMAVGdpdfvMrR7zLpSB20wnfxbZ45x48JPBUzZzVD
/CfQ5HjcdMOYcnjWFQ93VoiuC8LZ1I7D0h2du9NhcEovVxV3Ps224b0iIiNtZr4CHoo9aDtAljAI
BgQXIN3kJyGCo6bEz0gODTvgHUryZ2wm3hqj90eR32HHNHQz6zrmkHNl4CJ6asOCM5MHi6b1a+FU
JVwRSOCVY45c7zVye8lg2Q7AoMEa9ECKmIGbMWsEuY/MtkZ6aDD39ieBorA8TwoLVfXfYGSqvuEu
1jsCbhJexBfjtcSXhkMvHvPVTxSHuojBxUJwbLN4rgGx2u/H9g7sYtQP59EfY7suEFZ2z9wmVobT
wTfYNtvyVcekCqCXhlzLsWVdBu8t/9dagg3jBghg6TCtjeJsQ63AvKY6jrotcqq5XpOPIGqPYEkR
hKtzC77fwtQF+SHWJmFMw1kNvveWaJrxadSqAI8vwYKspuYDzCFyIfolHsNBDNhlicS/zgpmuFv+
vJeCQzNMYJwtpL+vJIoui8U2dAmr3LEVvYaoAg1aCNTyBXUMCoiSoDGQDDc7oV0fswQG5aFcJ6u5
wwshISabPel8SjPx14jciKz3SOQW7pkHDe5Gg9xJufe982Rt323dt81TjwqfL32symdXz8Ai4etr
2o+6hCt/ZXMoP3x/WhjeJyUp/Pn6ID7YG9UTRcIOM+iNRnOotKw3UanG4S4zd7omcJG/urY3tHdq
/OqV4d4plnzg00yWpG2q/QO9oG/oVocHslurAJZF73mdG1DMIQelSRnoVTkykJpSuCxIE83cyVsJ
GH91LiGuKR6CZYj/t6cRGALxiFfIulu36NXFr6FaT10GCN43Im6jytc9Dt83J9D6wc5syTnC0cyV
IOnFaElkDHyYKUMGi4Y6d9kiCNV2MQTezNWJvgmVO8J5KrSqW7nWnWiwGmJdBIUoggGOzVWpaNtd
8Gb/i4s5Rzm+4OkwznAeHKOyq1kZHQHWTzVOqbaph28o7dIrIG4zIWhZ7gVCnVoGc1P17satsJqp
xYdnfFhbtCMnx1DAEf/IvYh/p9eKo2EPaaYsBRW1Tha2/61z+sm5o1Shb0OE3eL2oBK6+IFF/t+Q
gCiK/HI/osBHQBLrv9KS1DX7zoWzWXgkR6fk2q2fyyxES77pJE0R8Zem9pg5/+9Xw3TT1AfxuQan
yd7P/q+tJHqfRpcH+jxoygAVkguRa5p/rUSXfpNmAwpmC05m8YfmSp/mm2CTJDV+Ff2ajI4Gayqm
rhpt2vJXcVkaiCEM+jjVrBFnu/jgJhrkdXiS8TVHmn3yTR5BS1I5RrqNdHquG2i9dsnV+cxg74Tl
uFdfLaEDri1Q8FO5KRkcoxBbxvx6t0DpNLGxLcOd/RdatOS0KxAl5LOg6SXL81sHEFTw3eVc9ilN
lEDF7pmH8uQ6I0LYXkVeprQnLtTfR0K75iKH4rei40M/VpxjNVYZyk6ltYAvGQPHVwkNSnK+vb6t
9EDviMr/YGmaEpZa+NoyI2oa5JnsoApq6KZf1ecpHT4LISoWJ8rkrjofYd4i76ceEdvTNI6qQ5aj
0lT7AC62OGGSs3UiMOYUHXKevUmpR9C1f1gINEV5DHtdBEfVzWCvtXg9f4bDx5Hvc9YOD2OTl1Zl
4BR7bY8dI2kUMFZopJJxDl+FRysDfxujnUW5hmN7CPaUIR2KT81M/lycNEyu9izL0UqrzaogfL0I
UBI+g0/k2WPn7LfGgerh4SuNJW1CtgKdQiIIWCgRlYXscu6q7+E6hKWYWCrgnmz1fWJPXws0rwRf
qNrGlVQLWk/6OTvd8HNMaY0uih+JIoBFpUHJhSICuHFk4zQmcM0VAntIrTu58dHSjLrvDffy86xw
bZcHCyR8xv4QJhQYWs3SvY7aDzLTZn+h0De3VLc7r1cFOHJ0wzUeJ/3+9n6SyWlXNjkHLCgiy8A8
ACN+N7RqnKHOM+jXFSe9ELEH6dX5R2Glgk8RG6tHbqlYYItxJuGH4ExkSFy5DzRylPaFxtwjfngw
VfJXVumj7vL7VZNgJEg07h6aRXYXkHRa2f0qjTxQq9Tvcf33OvEYUxWl2i/Hay37MoBWFjMlq458
7mykGDy3DTw3hKfCzUR/lKWxPMvy9MTFTqR2hWS/5suqgaC3z6kV10sBIba/lIUy0wkRj4bQiYOp
yzPtY2Jd1UAuaPM557ZKt1mQpdZHV4Z/j2dUFOVQ/0zl4WB0WYXj/VeqctIGJIJA/xqu3RF4HF8c
BcYIlRYJslInEz5eQZmbLonTqgW10YyLUKef9ymQKBJlr+ktoZ2bihHfLQmh6mqYJnjcw/sj0Vgo
s1Uy2oJedCNVmWt2jD5YgheEihSuEmUExlD+5cgTtp79Gw4gF9778eD+IHL7QfDLRVBV33BhjbJZ
Y1yVtS78k37HqcP5sZJ9oP+iDV/lF05M7XPhcrxrqUUNScZPg6NnABnVgXKAIiCBuzPqqO96F307
LdqZeE+BUHP04/lutm6S1m65++2R8w0fSnDrFZe4nrv8zbpMz32H52IvTYTskbGk/yjcRDR26gjJ
u9jfJuQ46FFIJEeEXYZIej2YTwzIVcFMMIPc0Pf+BJoFDBWDurajnxlu61k2t6N641fc1Iy4qUlX
9lsrVagTrBk+AjgcVTygXGdUMNqTwK4ahzRP01/0EeZTz1Pyl55CpQcEkl83HCswQZFPObQmKuyJ
Zm63BJVtO23VZvq7whL3LVqqeoQEBlraKY9lpsNaKbGRWiSf67tq/gMSSwQAXlmxDVxrUIAl4Ujz
JFsEMgIyrpnz/CVMHC+K/8vcUfaTHxZha/j7+sM8DZwtr6p7JG/xqZ7nUlZ817FXEvsFyo4+BtQw
Iry0uq6kEfLOuTcPV36XUoXTrN7/owEGj9I60zptHmnl49wng09uZaP7vwxMCntILZ0oT2ReiXhP
pp5S5aUIdLnVSuSBQ6Io0p3OjTHNy3kD+opQliIUqcsOST34JLnL64LVsGCbwSS5PFYVAWdAsa2J
8HlumV6fZrX3WVyA5tJjokyXQmRgSF4aKdnCV1WBG6LEGt09hT2v27PdouVj94NqA1QhpB9ONqoO
Rm4bIQDGUefDc0ssvsmE5ukRiGAlTALzBlJKFwdnsAe5z3Am6b/3lL/cQ2eqBL1Tnq+wTunzLWce
82X9uwH/OZ93VFqspryqHIq/ZXav1Id4MCWUvy4rnwfjRYJ0ahTswINCIKONwIiYd/aa+hsyjjOT
yDNs2A/8isbOJ7gK7kt2R3zClCrLCSKOC/Jvzo9lAtdWlNFVz5HrQrdZrWKvMi+VxEwXfSEMzvvm
C0DID5zMEnQPXpEF2NKCuB3a+HDXvxHh50/JA+SoE/ADZjtKm8UVWB84NlkJa+L2YKU56UqVtsik
DPWsmP9L9Tk5QEPEMYVPIihC+7XEToBQmsh5TxyAYUeLirVsgTBDNW3CwvQVCAOCYbAHuX8oqaBx
fjhQCYzXyTYSvBRBN/R08jh7RE5Zs8RsAhCyxmu73Q0/sjux420oDYzTgecv7Fak+5A647IAdxiX
4F42KdMtmetxDOawpQhr0yRt/tNCIw9IpvWrnxMKSnGkC7jpSX1dbKxvlZO2IOjH4i+qVspzOKXB
CHuHvpH/xjHQZ7eshpdrWFMK51v0+A5wuB0QxuHU3iNJUUxCtEEVgXnUxGMEOA9uEvp9LQbBkZSv
5jR97cucTL0KPfhHQVyfgwzIXGE3BZeHLdO6ScIOO8Z2pNg8ZJf70Wf8R/0dfUciW4/UF7nAT/0/
OUg3BjrFESd8tYN6o1w/GEt8MIcsuNZ5Rrw1XN6iULeuyAi5sym6x2E9MbD6CcYJG45XNB9z6hR1
R3mUmhjQUD7BqrbNxbBno+kaTE+Phvi2yk5gaD4ehEFNeFTajwgSicy165E0Qog3yXS/9uyYz/fu
dm3KC4PAUUdvG8QFjECKhHN/71QkR41/szAvNZ0QyKJ5DnKo8W/yHDh20pPCKOtXbiLJY+Z5NByx
qD2QWeIz+udpCM0cjAZg++FlhwCHBLSAumn/XPrLaV2wqKiJiX5wFcABp2qbtC4+GlryfxqFd2Y/
PqmN/uOgtPLUvif5GgAX1td8eQxRFP2Lx9ZmRMnB1a04IaURefkyVXH/3fa+1WZ9gAkUjTLMvmIX
mRjP3SEseXtbbiiwSeQHNqzUsUlUdfbDegqN3dF0djY2xFHN8gegDSlqsDmjUWpLB4g/Pqq+xJYn
eO3q71VKpJ72ZOYBjLB+muK0JQqz2psyGdbedMu67Qva6s1HMowZp8o9iuXjK/qu3K9FCIElAOnX
uAcFXLpWPaomV6GdvEycnYe/1paIaQS2weUeTWlw5uGn542iPIOd9HAplIArNLawe4Cba5i3i2wZ
zgN/A9eL+4BWE/83dh3+y62pnCwB0MN1jAkKOC4oEM66BUHID9S00t8tE6gMRjHFZkTSE/jVO0G3
kowvPDtqlYMkOJC0A21m6CVkbCblgLyqbvmQjoQ2bb93CPTMVwKIMcrjGCPN5XEcPw7vY4Y+Hm0c
K285RmLGtFbYjDdK+w+CNTXU7L8nyTRxJsx/O6vYO/b3Vig2JFbIEfwSG0YOd6K7D2poTEEMW04o
zc1Dcwm3TqUWxmVPRBSLTZkZDmDjOD7Wt3Q81BKJ4hPupHm0buYGOL4ClCKi4+LQ4r2ZYbNLWGDI
frSN5IF6bD0HVYaDOnXcM6xWdWKBgU/hRKxk8c+ntoMSr8tKL53AMRCQVzUZnZKXhl9uvzHG6Pn1
P+7uzsEIT+55Bs3/Wp26lX23wrL5KiNq5tZqU5I5qTYMCqEIzKL3Dck7y5mJeHOtyaRLPFKgMI2+
bhiqxBczZUkZfAjkWan4PKWP1oGSxCIlVRjx6XQhn3TqJfsWBPEfVBtgTO5//UNQRwAL4tCtFFH6
ce4nqudDr27vfXXNEbpNIh+HRFrWbxPPMnZhdQm4VjdZ+I4y+41WYaYFnxirAnTatBUPC6N/eaUK
Ss3XPlmyR1abkkwU82ErZt2VogrG7RXQtqufoIpk6tn3fzlnyx8tP7yaUek5L4y94TPpnt+EuTeK
rlB17wSqg3D6Ts3pLFVa2k0B7mdRMYAsGwZLRUwVipi5U1wZLJ3Y/tKGv0kq3+lqXT/oVWWD1g54
p4buBcHFM1v/yaImTcdSSKT+Klq1ZYeDVFm99qypSwgMEyx6Kgn+xEVQveu8XmhQI4wbfTcapCan
ydbpUoB/qAef3EYQiZJ+81Ax6OFu16MinmLhRnKLEIW6ID/TtsSPWdgDacrai+PAMSErvtxpb3n8
FX6n0NLp8/afkCYDWftz4yEL0cfO4/QRL09nimauwThWE5GqoxAvj84pQeGy8CCUb1ONLCquKMlt
n6MNZITSdUp+z0sYjMcC5d0VnHoypazXlHQN90aSaj3/9hV6Hae3f/rHKqcgImj0bLXUZ08NLHZj
r1b0cCcQ91wz+zsrP/PIpTgJf05lJOEoAEKNeU8AFLk8195c4VBvpSPvpfXjdnB8GoWjY9tNkwYg
vTnCxM8qmGvqcI7Fig+DBXsKqAPxAn2tizQuhoETCy38QVbB7UocP6IeeBO9UDhDKZ5MxHWfie+W
npVri+uSPYneiZbIrsA+bOk22GHnkP6kqbLsm8ZR7Oj4FiRgb6444RV0JdH7O2+m6Nyzea2o1QPg
6Jegfno1F8NXkWiaIaU0gjppL44gBKQBr57Y4XWyMfsIuO5XLR5H4bmS+77qmSgWj6XVJvojJJTX
PVD2r+OUCXD2aG51l6J77u87S5RsRwvsmp4CEPBXslLY8Y6pzIUUhgBh1gW7zy52cE++VzbDSS6k
SQ0hFTHEy+MMLwA3u8ZfN1BHeLXsdphP9v2dgZ40QbKcD/xBzOYlX8e0ZQk9etF5K8d6aJv2R5OD
w8VqvZkuMnNP6bsaYI51tyXHJUechXA7fS4Z24lh4V9S1JCKuPPxeHmO8yMPMTkWONXrcUe2H9h+
Pp+nD/M0heVIDv5gAKBOKiTOhFUopNvZ2QvBm6AcItbN1xS4OKH7TABSNkWQG61Vt5WqY9HDNM0Y
n7cWTo9CW/K3JZrJR3wKOtjHgUekvNKCQ8DFviQdrAhLdMbkBPtbAo3IbOxhKRHHpJISw2HjPXDV
3EVNcW7SSL+rjfrwZngwKUnUHJ0Aryww/cZf8rIUaMv0h4wvipwMsNG+FoVQuqTIzIFDYTLnLHg6
xE/s35VPpJM/W7EaESsnhqXOwZlJo2d9kEtFnbECfEuBF3XvOTi+j8qFbupirIoSYY/Qgv94+lse
MiKL9EA34r143g7Q814SBCDYYEtKk3lND+lPJFkidLPfnE9MYe5LlKZqv0e7R8iQzXZMKCg4duQT
c69RReRyYhbQOYZWQVrbmGcPks933Tt4nfI9+kPg1fqZa4oUwoscD/GsVa71tPm3/TuIY32AWaIP
r9gNnpcktp2xLPT5PBB0j4JAQCHp3705D+5Q7kR1VWg6NlEMP+sHWxcK94j4Cig9AHkalu//kV2K
ZuMSAD/PWd+moLN712AUEpJurxFEyedyfk8gR3iMZNnt4Rjj8dil2hoLx3yOUu7Ag3ZB8xMSwkj6
vE1C9ahX0m/j0YkX2scMSX6zhSdr0RRFvEXAvgMK70DCi7WLBQDwau5sNHyDw2DnhGrdLtC7iK+u
t0AK5alnNjb1dFBwpDgYuJETTi5Jbb09bl0gx//wskfrexqdGHTkcCWrnVFt+Lfzvk8sOIzj0hmg
7TJlxs9HeepNDcj8+9eRHx/5UAs4rKWsCjBsyI9xuYpYI1aoidxc8QZgBToiCRG/Gh5h8WNrSFZu
JvBGPu3upLdBlpqS+13qO2EdBbbIEXhq6dQd6UPS1ePAcZ6xhkwjebFCDyTVjviEqq0dbiWsZjqT
rgTdl4fsyj2V4VM/lItDJKHpAvkaMlLqf1W06QyrV0kNpKCwV4jJ3JB+bX/vBsK/idlO0LyeaNuy
/GSwUPn8g1hnMCt5/nBgurpe3ainPUONDMu9PKZ1rLINuOG8QpCRXBQuPMFYfalC/odvs24XUNts
EPfUoWWrqZGzS3N6EhdW7fw8jKKzT6CC+RMgdLL+FIUD0Q0aY7JUGboicPo+Wu64KHPeCChqXBoZ
qW04+k1gGkCueJSk7qxtZtla0J05jJMhQwgBWjJLzrJvuKKxYbBCkuFGUxWCSaEi5QiGALhRYrLZ
+oqyqih3+CBniQ3jBL13SSr7ZFNJFruG/P71niR5dkWAnxY1rWDDVb1nEtLNd1mid19REmnxusEq
afQkZoyqGE/4W9hayp+5mnrxJ+dx5UPvVseuwXip+7aWHeTAxbBe0YgcBBv9t9BERy7wqui7VC6/
vVJOpQlCwiC3XEVZZrw8atBvxCF4EtIWOGSHns9L3Vn3ni/9U+cNTtSH8W/mP9n99PdT4oIXDtcj
Kn7Rr79TiSZ0Iw3xisygNWaAroGcyr8r4eX6gEXopt8H6ZwdrgkN6Va/Lpa7Z9xN6s7GY+CfLA4f
XXI2vaXKfnFi5xxjuA9yhlxCEQxfOBsX6MJ9ix4+XeCZWd7AoHB8+7nsVQsniCy+XO4QdXLFpgTd
I07A8XFLkvBA8ydMyWNYnlZILiUqLPZIi56loO7yJHu0jp4JcHVRUmd6CiiBSXrVrJvgpdA6jO+M
Lx/5qfpkEFiU6SzGvhvlDbROn39uBxltGCaMPFvD5eZbHzw8YQHoD9UmllIAe9g/L5hgPBuW7B1I
u9vUCgikVwKUSNFyuvLH73qc8q+RjvHmw13pmeaair4WQ5hC3JptJ+dqY/QtFHyOo550CMyy1ELM
BpuIttoT1A6V8H21MJEuqsP9iM45azXbZMEkMnNcy9x70eynjmYWUsFMlk52UApEfwcyPfzSK2GB
oUzdOsBYJbWPTJbNCGYxTCxadQswHv518hYtDVFC+eHeAEAeqMH6GeEkNSSG42B1sJfcUvX94dAg
o4+ditUgAMMvwQgcaEh0sA1julMR1L66SkIXkMWmN7AqZXLSW85UbrIUqoPwoYLwDH79QbvvpSSV
xYGLacWMqOoKZxMjZV90+wQh1INGmUTAvo/IKYNP9zPly5KA6KI1fsFpI9pvadjiRL3NGSQDIWq3
mP48dc3KYc8PDcPRloBX1wpV3dLSAmd8WHuuYy823wBW/E3ZAiQqQIC/vREVKCyVVXcT2Js/IjZu
le+yvPdSjuQdgBktwwzTgh43TI0PizCAVmv0xy0tbUifzk/nPgPIcUZ6grSLx8BisypHCwo1tm8V
nZeGAm/vA/ZWYmxYDp2ZR2544bwbqvu/B/x+tMfIUy+kf6627W0UZnXl9si3wNHouz2GG2UfEAX3
nUsHk9phTX89gadY4IdiWfQUt0sZHO47EH+N5u3LLXzePPoRosMMMv4XjI28JoH1BSzgRgdkEt1a
2rp9d13O+QSJ7prE842lnSKqde8LN4ji1G0PDN37xqd8UaV35ege1ruIrY8glqqVPI41TjmZwMWA
W73t1CLpKP8Ion+N756Ke9WL7xei8yHyFDZRV8fnCprNy+CmBB2oABPrEjPeqIj4p+uxN1xwwYWe
GbnITjeAzSVUgZg7pxSb5ZmDxmAOJI9Ju1sw7xgpLhIFiE4wPUg8hMMSCPMFeIsls8cbhbEu5aJ6
s4+kYjjtge4Ux9TyCPnAKmTTFYcHL5Gy0Vtu/O9ZQmBn+Np/1nI63Q/ekPNnBjsfalFxDmQvo9Sm
pa4SPqb4TyGorP7nsbiL72VUiI+9j4H3gSOAtmiVoX2eIT1/ehewCPoEDG+yEyxengwE2qZID0bq
adjOlbpZY1WuSPqEhkxZwWHnrLw4lmEdO7L0cFpdKuUMGZghr/+ve91jUIyEu+YFRurIQTIG3qwP
GTACcGZLkwjwz6/9LtFbVzKh1VhIX8s0EqNsV+mqh5nO9YG5LVaJvx9HSNRg2XcIQmh27aln+5zG
ZQnVT3pjkzOAKagHn2WumqTu9MiRPkDPQJbrFPyBhCWuiz196BVDqU4wD8+XFDn6Dg1q3SmBvyYi
BVpeDH1FTqozbkjEB3zJruy6DbBWbNmGi+gpZW9GgUfeZFht6ApAE69zOLxQbZ72XDmBdBII/5Ua
7r6rxgEZCcYRKUqFeide6fDJgpQ9IotbvOOCMjT10Tm4AABOaMkzrSlPPaLnadtHKHjsysP5Z7Ky
a9drzEUl4IJGsqeIU1ug09lakKlYtkjTMXg66gfzmiwyVqwQdsWgSo86uupHwPXaIOStnhFQ2TYV
ZLnxggMLIuIMzkRTLK8MRjcwzXLkX8K/7w36KNT4iDRv/LtJ64kx86GejmtYoNH0Htpx8nzHMw+n
YfyTx4XmhAnDf1Yy1lY8eM9b2sPC1Ld8oSPD7RBd13lnJdYa9NHQrUeypvF3jMv1HFSHenlU6g4m
daVziFCFR0+eWJoS3M7e4r4kNySxnRXt3VwJtSdciSlbLrZxRG3cUumYy/7vyuwC+iW9p9rgIK71
sOgeFgI10NpGlLFoLBalqQIRxvwIaRHoAXYCV4g0LP02dRT7ViarGPtsYU2UGI+wM4beIKY8fy49
TxTs9dT+ioLcsNlchbmYJDuquA0HxhGojpAVtwBnMAnOR4xyjfLj9T9phWORhoSQTE036o8bvUnu
RUjIXefSfNjW5sSh+T5o2tLgh8lcYOd6Vb+9uChf/QrLv61FXg9BB6/3AigPCqYdIYgBxfRPEBwc
Fb3zdKyTlcVXa9orsrDn+QC+Khsg2rVjDH6TbQen4x6BEW/XCi9LqCYMfNm8dGW5y2PfXKzgqohs
1ZUNMbqV3+7go9ShyDNu1OylxqV69UbDtUPwhppMfO3IDJ+USpngvQOHlwKDcsngX9DZm6qIeNhG
embyx1Wt9fmdpbi1vcru/LnXHDpEcc3Gyqnkpur6mwdKucas+1fcQc3G663WtZS9HoqhHPdqjgR1
j3PtMyTbCPssndd2vgutt1dcQZefw/ClqLNxRg2ZQ1w0dy1DulU3rlSK1gWBKLBPBxF3nbLhoT/v
VScH/w9DaRtkZZO3u78ekDDPC9Ov8yR09JcUdUI3VVfAy3DTZXS6znJ31554xlyUQxMt+G2HrPef
omAPengsjFmKvWA4OXhfAQ9jBpUrf2ap/vzBkLMH2XMfo6gcLPZMi6vMJvaZl77RvGSQ1JDU57Mp
912tVsyhxMuMFO0ux6BhPoHNMm6oR3uR4uVnFg5ZNUKAcIv3Nbuc3hU0xnNiP9FswBu+/9iK/Pp6
kbclwRCVBL7gvX2OQkH+coTAhYPwB0hmw90Qrg1UBuHqOZv91Frf87l7VQZfG0qxf5b4sgFz7fh9
48U9gQNkOHypyYCd1ZH8H8V3gnSPf+xrUdeNzHems2A3Oq2t6Kfwd9FzWG3r5PCmORCw/RxDC3Uq
37F9qPwlOgsdgXbVQhXNnS7eYrX0OI1bHjfd6Vm01l448CZ3vRcyFlj8e1y2+pSuEih7QYKOyFi1
M6FL2UUFpef/BtXoZlsPTKYb98GJx0tQG0Y5uMWW4m/H5DC5/dkSgsl1+bTcF16P4DOQMKHVn33b
x74XtjhjtkkdwygnQO20M7NWotnNGqPREfibF0uS2e9K496vwbZ+YWHUy76Zt/G7ykX85fQDNCcQ
FVwXShTf1BbzMP1RdQF6DkaLYiDHJRsda7kg6iZyqLX/UOYVm9SjuYJe2kSh0WhKNWRbvB9fuIUa
aTNpU+tm+uh/8DClIObcmoITENJbnus1K6nnP6JvjhnZ60+wFgYkFfQPjRfEoCFWbXlpyDZAWvoB
IR8CQnXNHQDkSm9dRyqESOXTwvHdR2Th8B3mU+fVYydYWu/M+DSMVP3XVv4BzcTPVZdiZnibECMD
QfjfgKCQHJC3GTruExOzcqN3pjeH6Ch8GoP1QRPkZj6bmx5lScy+79ZfSn9dUPnjoRsHR5Bb6t+n
cOcI7LNYkqroA5obHBL5En3w/Da11sYRqEWnEdBFri6X8/WDdA39wCSEevPEghYIPx8362wYEbhO
4eUF2hg5bY4SsZ1hIfHaJg4Blo27JDu9+e8EE4lSRgP6qMub2ErU0aZ9krAsAGs4pFW1PZ0Y+pyo
kEAtr9E/qfaSsXhc66OwfZd7Kzm2HNQOC76v/kv6EKKcjGxPokLDMTm0qxaquZvmWREUmqUhuqHf
eF+gfLymF5yzU/+89rCill6N4vQdy++6itOVntF8WeY84YwSARkgDVqXmgj1TOrfPjg/8XbsGbDz
f49TRprzjqRoxrPatOPQqnoVraOcpG7S3daZaz05CD4a1Vb63T4mO8m/wGYm8E57TiQwrgmkk26j
79O3L6ObPRhZCos1jdTwVLIZt++p0DaueJsmzBk6DqaN+7otme2BcYRw/KcnDtX00N5BPXcYaC3g
nO5VCCt/gApoS5CNR3HgZArSLLyjjquagWB7jxtsNOoScKNnJpUYmSmc1ZNiKDaV6e1I2GgjA1OC
pyL5ytvc7sAwepiqxt3qRdz/Wkc2o2WyXmyGqxqapVqlIR/7NS+pYWwoWgcEXyrtNT8/UzYDmymB
X2TlpR/HJ5jKHehpuuWdOccN1burMLwM6ieEe2xjIGpK7s2U3kUO+Zjc1Wj9BW3TREfeVjGFE3jQ
wVvOUUIzHdCTUrUY5pNbc6BvZWJiJvuuRdysSskYgE5mXquCw7esfwe4Qvj60ai/q27OugZBMOvk
e0nmw5BQ8YVq5uLZU1F3WyivuJOBEBR3IEkU7Kw9uCJKLwAvkewMm6rPPLq08368Jl53kC20Mc13
pNeePZbM11FSv5f2v94OdEUj5rYOdGMnHiajlP1ZobWIYqLt74CEiJnyeUGbMw768K4YCfKIGC/v
cXQep/O48aUIW5QwRUSzqzCzGWI35Ib6Xh6uEivL3O9dk5NCvGFkXf3okb3Pgi9QuwYSmnM3+pdk
kP/35QOuC00RXQRD/h9ubKXAhAB6IjyU4p8VoYzI+9Y1/mbouJhADbj3qOYHCAqxZ2kUx6TQ0Ofn
IaGaN7NajYYquadTdaXODwWcN+/DZ/yCwr84uCOpSOo47Nm7bfr6W4tOgDyA6c4DvN4BFne1c7Cj
7digW2ext2dVmXiSVDZMUtwg9T83Ar/fMNjV68OOA8acytEhTf7XgTHJMNpuOv/MibkRfo72ybES
+7ND6jsl5E06k7TnhFYJpVEfO6YFcderj4jgiPW5wExZKs6N/W+Y7QsXf/eI0ynlxZW6HK33R+G3
prYb8KJbzUEiM1rwi0yATLnsj+naUYV7xBnDS2/N6+KvW+eja4wbU2MD/b5UaZ1hJEttdr8rOivh
IoIjqJ5YS/S4kKe0WkzjFsRHcYHe2XG7bm8jWWjN930DcuYYn/5w+Cu0yml/Q2LbyOHcRRHX7UNx
2vfkgfQAOmAvxLeIS5qtnklOaNPJUGfD26C+Vlwd3eL0Bh9tUyuIhFicophUH6NWupCpdygzvTLp
FYo6gpBt5+o8mP+9i/XkIIKadt27VCllcZgC+IVLEuAh9D4/m+YFS7zgfQElms6A7+ZSDngCnV80
3ZaVp+cooc8OmNO8U/fJPJ59o0QXq+gtvUUpmRZpniInoQpkhJqHoL7LIJ9RFI7Fobvc6nBAcsvb
BOvALLG1pSfvEN5o3TsHVBDz7SIvD4pKfVImLE9rEGyO5DEN4Vj/E4lNfBax5Z44A0U+aZC+GGjo
F1hBoWGUPSJ4Yumj+AjdxrQHqQSeWL9zMoxplCzdzANjaVw3UUpK/w/qC6QVLCcFjFGxFPSJcU3L
b67R9Vk5jOoQj6wRNbYggcEs5ZSR2B+DVCPgO4ZVidRkSlccYRD5FFyh6dqzwAYRJIT5f9CNecji
AX9ZN819gmqaW1wYYiR5Phbmt1UvzhvLVBnrNbJp5tJKRDNZdtMbzXI1FXMDI/XIiFQH3slq1XvV
QB82L/UvGd1Wl3QxnWF8/n1nTng1lSfmRmN4c0qn5YpetmYtecIUPh2A9grs9UmYWwPpufB/npyt
xNwY+/YUYX2rQquWTSVOxeEVtqvE53Hd8PGDUMs8GKlUqWTrG6ZTtdR15jWVtTa+9Q01z/nSvmba
U13pwp9C6omZzQlcUz7VFwwOCOfJJDdp1/hxuBQBgwpZcXGZ3CHsBMew5zvVUJmgjNQ65FqGNHLE
kybR1S6NEINszauv9AgzsqJN1Mb+v+xw2eol78wImeO4KjZAMcHWjw3Tkerw9nQrbkU0WbXvA8qO
jZ0sAAEG5g4TR2aFGG1FMUHUijK1cvaDrQ5JrSKtXIfsngqEOgyzQXLv8bXSiz+tg69PTOwvkIxG
ZmNiFx4/Wt1Cdd8kY4YMkhncZulZIjutCT+Ha69jkAT6g4CHQQ68SUCOvUo3DwE53te0MWUSBfqc
QCDCy9l9/3cTmAqmnWlie+Gb1+xfdDaFnNk7EyfCIzE6kuI06W3rKD8E1szPNGjIiYWmnskGbOtH
Vp6+Ry0QnaFy6eGaCqfVkhSY46tSbdJOCklKp20DWBMawXn/BKu8lR61w9K18/5o8+NPF+5OKHDS
ouIsTilD68/PcNK5jk3S1QRwnioVEg8NSYOH5R2O1W5ru9uh4ieWS+dhVYkCVVU/keNs2KoQAARN
BrBhRrNBX6zVL7ctO906GAdZma7finZLbWGE4+SlqOKb8JBgZ5T3Um0fGAtj1A0A0/RDAIIAaXTB
Wf378/ucpCgL//dVqbut3wFRmyAT/oaHyniHTERFo2xMi6sqWwRYvpdHLFBxt5fCGujJB6vfK7if
c+YB2fPKUiArCTE8T53iGa1vt2bRqVAgFtoVINBXzP3falALkfVJPcKr7XWNwKSkMWX5fVyUaRuV
YbsFzYEa7cVWDZG4XFhjR+fHZWsveNb7HDhsgolbq99FZJpMz+hohrZ2skuhhZgSyDNnrNKPWzny
4D1LX01dhsaIaI/lmMJHYGDQKaao8FiR/lh7ci1U4xH0Y9SKVH1PDUMzMnUVOFktuL/k52CoIAEn
nWhrZK1/bhqRWznPeMGQhP/cmt/UclfVSGozes7ijE688N9l5ax0wSeI1vQ7FJQUTeLx3QOxtnxk
xXCOGRB3pfOUYQ3t6TCEfjrSD74Btg575Qu8tKst0ryexYf9Z/X50MRsKACqpPqLdkm+ICXsZ0IH
YQvAAWZPEEXdDrqygtxJs88vbGDWKeIaI97Ei7Vzo7cwR4IJKQToWVcRO8jxt3V4p0opjcbBZDRb
rXl/3E+3pXfSSNgPzG8RTHNRJUdQmS8gNnn6+716sTLeI0BPbXV/k9SrvX+xYidNMZzsu4HTU6Ia
uAozUyYvxK1GmGXIV1SFiv0sauzs/DWquMMs1yX4Ly6L1vM72zZDK61glLMTB4Cz2qFnIoISPdC2
UXvbW0mj07dMdpk1YgTzOJMX+C1MBKQurP03y+oVH7nP+YXHuMs7QwazlyOSNeEGDPnyn9uWsAAY
yI8IO39H76V6UDokkaQ8dQyFjbgU/90AYcdmipqjo82XfR3j8hziL0LCQEUoJNkqNVE6Te92R6CI
Sj19BOk3JilizvcYjeDA2U9L8pp0qk6HbXVAhEu6wd22y8/0G81BGTnLtNfd62tMvbqg2PZAD5Tl
Szx81fw5PUNcrg3xH4VGNce7sXEeeqipABso8l2gG0mD+fqKGwgAyYw4LMzWQgF8kq5TvVtF0sLr
ez7OYXHaVIJBQbcdIWeRzZz+YmFJJ0OYzZ9/5ZDxAb6lRrNvK0kSie3QbHC/esCcdnhYBQijXKNr
SSL68xC29ljsB09o9kdIYHCLVISJ8XszBPJKJpeO5fvEEZw2WezxrJSkAJjVCdyp1XGYy8yIE3ky
8+8GFKs9F5zhySCQ9tTb2DmVpYy2hAi/srPV5jTay3/64+CwRM4QKWa3SadtbLm902smAycLk/+W
Kk+zqbmgU2aIgIkoS+g1AKAcBBGeBm6HwaOn837Ce8sUjVMN7W1hA/Fwzd/tia9qfM120v572pa5
M3sf402WB2yrE/ciHIHTiVhxzURYmSL6wC4A/gL3nmFVxzWhWxBRm8ohetUs42lh21153/4x0arF
pX2XDZ2pRTPjoDQlyyzIhnK9XaMvOyOvCkeK9oHYjRQgM21IcripKX2fcGWh/ItHlplags0xclTc
VzMxB61MNjDaupGLL8hE3ZU4zEH0HmAGLSZjvpGdV3JVV2EgDEzP2jDfaqJWYZ0nUpFZQuK1H7qh
iwWHr25FaFWle/gTfG8fAD4Bi/+bXmCULmBZwERABlfheITB64nw0ySzcCK1Lwl67QC+BNSg0Fnm
2wlpQMWjcRCB/xGzFJ0kfnzqpFEvi3mgfKWo044LAcK9brGonJlbGbJdz/Ty5QJSV9vCyRV/fAgZ
h+r0geY/HF9h3FDKcrRTXRgjglvcRsbm4DN2jQMUIOjTQ6q/5WKKIV8GWTTYCAphonWHTFGs2TP7
AV1ODNvKYg/0oFrns3r4H2frrUJhFqgJMEVLEvZqdFxbKVGbsSvdS2MePjYMIUeWobDORQN8pOHQ
OB4DEqh36UH+jANvD8JP0Gekh7in/bXdk9yO9vyoxuN9DVLdaFgsSsacP1VEqmzFH3rGUez5LkSA
OJ+xyCSZ/15VwFgYq6gEbH77q0zy6/DPzw8BtcYWq+EyoL2Qg1no3lHxMthzy/oAmcZ6JUO3fMT8
B0eXah0RlHlD8KNLgAbPdjgmxsbB3+xFkYzV5B7iQ4nUTzXtSUMXVND2T6M/9XlUiPFHZYVok4Ed
vlbVG8YXY0hvoB7PfNaK1Hua7iMyByqDDuXc9T0q+UOxkz6+kyZ/g1cvBN6F4bMCpoHkzu9aDo49
2DKpcO4uuZyB5DHfuhnP4D4rzomrRCphqztCApF7wcd3nnamruzPSxVSXYDcHdPpxYkdiyb6FiEy
nt81U//R5Rd1grM3NYfJxFYiJWyu8gRHIgKX7TN4qBMamOgNxQjrAWw+zeF/yfSQ7KRNnsk94ReE
hgekIyi3xAo7K5W4X/SsqnHjTNGmTw0Wt6A/egbhUohOkWIWBM8QehwCTZs3zdOf58QfRvNXY6qS
nbm6X51kXMpC2WwnpLeqr0sfi+wpHr6CU9oRDv5RvcZ0/jyrSwaAO7wB2i/Hw1Ryw6Gv3uqUKSpQ
i/siXl3FhzLzwXpCsneXwDXiMLm/HrJFWqdYNyipPG7c4ubBDXCZk3OBAE9UUHUSW+a79sssa4Ce
8gIGy5cMhmXGRsqOldtuzAfG0+XvzbgfP6aVy2WEVmmTAx3MnyxkDg39nDgzbxiV7PCVFibTu4b7
M4/5wxn+JMgcjPH2cwToRNEYNKrnOX4iVhIGOX633qrxyI37ccsxB45YRwqC+YEqGN7BkNUoMdTL
63eqOMMaa3DBD30A187IaH+euF+dxeUmlyhdPN9yA2MyIrDBqCaaetFVnc2Re5uiLJzwAHRpM4ig
Gti5pMhOvTYOAoSwZniLP1317oD1LTN5auU4UhcUuznK1KhKcDRCsHPkNaZKkFU+16eym9GrHH9q
K02SPqU3JUIXH1kLVcnolISd9s8XXNIB063uHy3GGW/dlDHDNnjkUMru/U14M70HLmPr1aNfex3L
O7KElQQkrUFHtUxMrnn56xJXwfrGQE5OZFsqeCw4/+j5j6+QEhoknmr59d1RN9MioNMUQJB5OY/y
13LS4F8qIwgZ79TbS9xHV8ehOu/uC3HkctusGQk5ZNEEix0NCUAFWU/CFZ6Zqz8r9cNd0U2m65JC
K9bsCmLqAYwdBEj6Kb5bedpG808Vfx3OB/UWdaBWUg7xU79Fx4sU7uxiGps0HCWF8m1X057ZVMXZ
65M5rtJEOlmCQBmqdHjiqxXvETRRZQ4lSLzZ6350PNEe5JymyM2si6oM6Pe9GFZM9W22QCM2jUvl
JRr/6hAYku+TaAaS9qzz0+RhS+YaPFk6rdSQ1u8JMblxxvbhUigCTGlkNXMWVHyav9k7GJ0T0PZd
eztdJ5wThBFdX92jtZZxT+5noI6lvprfy5uIgsH4KYC1spfD6UEXLgND4lGu8Ety1gSaJA8i80Tb
VqCfhVynNYAGJy//lpPkDJTcfYiMmNP1DLnKcK80CUUfyC1BqmgYHTPonu3zRdaCYHV8Mgo0lo/B
h6HD+neM5UFK3KUpw+0b7wnDizcVFwcut0vKfKacwQg0FfBuYwQCY0J9A2AhYVDFp9/lNGfIB9ps
8N4G3kCvflNHhKLVwgMUF7AlMTUHq/2FbWMM1Xsw2ARxs9WXyiJPhA+QlR9C+DmaVNllHbq2rxhz
ho5UVs36gdrKVR7piZU4UXZusWeWdVNQ0JU4NEh49v3L3FHiW8YlFwJUJL39nASr9yJrKcjCC9yO
czcbEsJRxplVMqT5CuaemLffSh9dLtnaDPY0F6ZdFIRVDPXAddAvtQr73ju0CmXjkAd9PiBibi42
QRCS++0zJU6ZDk9u+QHF8qdcBLMaBaAPydI6+R8yzf4FsUoqv7bwXEtLBY7xezhStywwFseDBb8+
fglXFvjmM/WUawsaimHuaxvfi9g1cgUtjqLIPNrzPqPvY6+w9IaVl6xqlwgeD5sApShy1OYfVEO0
ILNZVBRcO023tiqr5kNg/jAtZWQg1hXupGk9CEJ3VtEN9etqOyVR2TmH4Qi7fpawUpVm91QhSase
uk6R2lwzVmm/pNZWHCa/U7O8/joA6bSzF/tbbvV04IZiDjUMS+4ds2dMeBdiNFu8NLfGeiTPrqX+
9oaebfHMafmRBMCJ4Ge4cYpxYTncMZqRnSZdaxGxwVmf2h52NuldUg26YEgWUOCdu5bd5a5k8C3r
AbmcFup9C/+ppbO93MLECosYrG5UNm+STsqR4HyK4MUe84RwTY7fO9a/f+TyQxj1XOFH7apiOHc4
P37pyt4IadHmZbu5oRk3mTjl/m/uIwQtoMTxg2suCoDd4zpR3IEzzcqiCGt4pI8gxk0AKKhKJY1b
s6vcQAnoEirRcygUId/iwhzJTooYlJwpwfgUE0c1Jjua4rhdj9J2OD4axpn/PpykllYZTdBf3j9t
e4WjFfr3E814Y635oIpsbPe3svw084jHZ2n6Q55xIX5bIZB7iHeFXwz3L3V0KV6pE86OifV0tVpb
Zm8sPnqZp6XPyEvEefCeuWbP7cI75uamN/IE7r6gufLYXVGzV2v0U+/C/WidXTw833oAr6Ifoau2
joe2Mkb9ktr1xYXlpO+6/Wp/MRL9glM/GAat2m8zo2s65U0j3iQuHEmKQ3/6NcuXMU7RQbbhl7Ya
u2RN1Y69wYP2/tzZdi6bOAJry0kUWiE78Q2qO28tO2QrTw2RnG95NlXZNS/SVw5w2kI0UvjYLMW1
iRepPR2NZEF/1trwqkEy8ZzEpdA5Y0nZYgn85TmH0CcpBW5GJNZrMCjHJmxg6PyjA+fu7Rr5+bYI
gvFzEJtyMOuHLzrCpHS0dt+u53ynrwoz2kgpeX0q/1YEfrg5YpcdPwb/DpPvaTsnqZKHWMd8voga
XuwxuRYXJH5E3AfN5byGlehUxveikpe6KVwuY6i3OdRnJIegO+Znwq3JJzcyX6QamnzFxV7RmTH8
If27yRtVpL8A0zqBmlPwtTc+PZmiWcAqN80p5osOmYpVRFJTbObowtsGBWvRFx2tuYSlIOcnZZMg
3ns9qXn2B/oljZy4yt2LMvUbzLItX+AiRsdWP8Jcjr8nwNdQ3i5PE9xXGNgE2wmLeXWDhKdMpPpC
n0TFIpGsYg6O6kepG8d13TiKW320lfom906bthKW0Y/tR17E3WCwyW5A9/EbxZvzC+dbGh1bXkpB
giXSXj+vEUmQxrOWxYgClY2VCAFuOJ9qWQ7TDTfkYPe8vPqEEdeaEKWefUDCvMhos0KeEGB7yFHO
Uo5CLr7zJcITVhFXabDO7Vvcf53h8uzSFz1R6NZjU1KZOcs4GQ5bDbyrVuwp0tB9hRpknwtvRkaU
J2Ii7oV3PmL1IgUf7nsVK11FzRSgV/6nkvxlewgL0EG0ozQoJmIlMxA4WExwkDsYGXJfu8gnkg9e
0gJkKuzsmui27iW3H2GtdVrvGqwbBiZ8L5EN0qO0RM/XH0YSdnhhKLKt9pu1mSCGkGYgGdaFC0DB
zB4l4a5Sh6dOfo/tDB7fn/arR2+bFqTk1I2yZ05xfbUukL2lm6ihB4bePMLtfYx+A7/Vc4BVPnXa
/rEQc764SdupNHd6dQYl7+vyxm3aRESWXXD0ySGnBGaucaMJoDT3Smgp9mkuV6+yrwlVVL3kInnH
757oL/K/6atPbhWDQcZSCv20t+E7UWPYPGp0osE9NsYQul5/IinblgG6oA8hSd7hulZPA4teesX3
XImmyo84OfhiWdQM4nbkhllo+K61g09S0bLZa4sDeh2gpBngqFOhMeNzl+TgxNoWmhhHZVs9Hpi7
PiCPhlwTUSjNWgXQFUMaNtSnEwHah+EDLNCb/eCKXCpGW4u3EvlLjnZMev2ZT/C6Lt8px4BwlWWb
L8lRBrzr2Z8k3bv2GMa85YaWfezdnK3uclnW6pkFHubeH8f74Q0yAx/0FBuFQvQRgyUmHNQ3GOtm
fjUNeLtOu7peqCCsyJiKsuZo9phh7WE3wQF2kvkvfz/y4ZFaFSyIW0ADfTdMTbFk6eNqLZ3T8DSb
0GhoCsYZelffWrjDOLiut/f0cEtiKN1s+whiyPO+PtJqG7h2gB7CPrGF2hf/fcy/PpkyMzZXAWiH
Aq+ThfQHSykFSAPhR/Q5WsYXqRdKRbF6jHG2YtbkxaFC54ELwKlpAy5yGjwdwmQ41fqtpbRoZEpn
yiyhCVTKQ5AaMLCh1dc4AeIBPEnhPqLNE7+IbjE2/sOa63WCOOSW7BCtHm9RyJoNcqnLeFNkqL1k
NsFdtjGfzrVM7avA9unJg8F5OuGL88pkgPMCIgrU+YbvpF+AN4vnMWMdcQZCM0/omyjtbr4BAeZZ
J8BexjE/jfbtQTrMl7oxWDKKgOsPTrJGLv4/07ETZ8OMT6rXbVVIO4JiOADUfJBNvEZP31EUuu/F
IBMqhkYL5o3bFqJihsrEHC6RsOqsFYmgaoQ1dhb6BpipjpVTJSxQXgPO60AYzHHpkGo2kKJT5nwG
pJJqgmDMixt2aidXRKnxUfGec2X93AxNeJiGDVeBiz6cE6bg1aVmMyDuakWi9dHGSoQ792RJ+qWr
ccbBdxjBVuHLJvVFsMcQE0a5+fyeW1GC4dDphgiXmcIrSl4fkkiO7Tp4zDTQgDhhORFf3uRzg8mx
Dg03CDyBSNg0Laj7JJ+DOrnBdrx47sQbJLs1dKtyU4dXucMgR/VI2bg5o0iOjgHHRqwgRNxi5C7P
GqvoUBqQki4hcHIhgR0I+dzqisz/73pOnJcVqGy/+cx944qqYe9mztIItQOOQrXAqoGcumJMxUib
CKsc1TYRgMC8ANw4V2HwevzD4u6h9BqbKyi1uj0KB7ScAbSrw7Juo+2GEssGakPbceqnOZSJq20F
ylaWZLKO1Fui2pNWcrz27J7EEV3cSCIdUt6/DnMoa9WxkW7kWpH0SvpFcPxHKsyJ9OwVlFUmfbxg
FMoimjpe5MGnnPAhWBZpdxQqcQPyXDmBl2DWDaPP56PBp2g9S8z5bzoGlNALW55NZqqS4KMf6jRG
0ROwIHDlWUJhP7tveaKp3YhcPwBnIcLMSG35y1EBRqtiMetIo71KN8ZnEtEyYI2bG6CAjOZYvbmw
sbIYSJb7FNdGc78LkaOaPuaXXtFq8YhLfIRBfKvKtomKZB5ZGKLi5EVm/YwSh/f8izBPlBRa+LV7
SFIbr/npFYY7J/1AgRO+3Qh6BwMEja1JgMqf0DvjikNn4+F+JR/VjL/vn2UDelA6l3Hpeef8JoBp
OYHqECtlexM8l9cFaMG7n+EHIOPQerNoGvZjzlo2GYqQtHIn1NfHbqVJCIQ8Md7A/Wap0v04Civ2
crxMbFSfSUQH8WltPf9lEPPeSVJJhSUHZeU4tE4DAAVUYfdsn0IL/Qx0PtQuwryxgmZRgV+qJH/A
bj3sA7tjdfkk17tbz9gnkeN73U6YTtoKySF5Pg/siPySfXbOYGDgV/56MOz0WGdMJ3LYzliqN45w
cAbFlGQ3RmYKMwT0DzWCOv3sGuiNWDou9Y13EX6YKU+jIKJ0wI08o9+Vc3813r6HmGqmWf8nYOqo
7gG/AF31BOnmCXgVj8DFg9ZT7IWQs1upKWSyy30YMcSGVzNj9L2/eNIdLHyxnaxXf53s/UHykvUp
ljETqm0N2vJJv+FZ7x9MtvK10uMkFQ1iATsDEIG1ZLYJvoT5420oKNW5jr7OPMq5p1JN30eQEvJ9
UpcbpAQCRpR8AUEgmH847JQqeBICvu3YT2qXd3pbg1uQR2tt2Wc4nxd9fTPr2bocVEtl7CeM9UbM
kd01Op3yIRC/mC07BYwrm34A/x7gGQ1p5SsB+8mhteMS68u4n7147MKPL2SVRSoCq1Wq0+MjKdfo
f0bdft6bvZK3dACgxsXLAkPcEIl1hansKeu/Tis3QAQ9TNiiZrPcnMQZ1sFrvlp5ARXe/XOBSynZ
BY4LcYqCNenN+E5baaZfAknF9Sqvs9mHWLCLi1oD2I60IpkpPj9DZWQf+th4ux4ic703sM03z7dH
3Ac/bjFY9+Oc+Yd8jVL4hniuTEcmsEnZKQkB5TxTMfGFXgWJQMb191FbFwSL9EmJlVqMO1DwP1Km
KHf8vMWwTin6du8S+AQBXeppPSdWn/bU0D80QMFaagXitUlOI9mP8lJvmpRvFA2ls5f32kPA7i+e
dWMyVzbtLuWpMTp78Y4WLg7ClQXAplQ9hN5Y4ZhgirejdIcLX2cnXIIjfhANdP/UCHL7ReK30jsM
9VF/+AosEDCzY75REg5LK210NNCASdT9XlP986FzcO/xPrhHWb3G4l8fyoJYFx6mk4bu0avRmerg
iZ2Df0NKayAKbV49G+OU758b0hs77Rcz0VFv0oVQIy/w5xHXHsk2zXeDwTYJKnVNKKCQ5Ze2BITO
expBHraFZJqjmetO0NF328G8PeiDYmO+yqLNOJJUx6EHduJ3y/Rw319BUumyyKYQipNezCF7HbYP
ppWpWJ4Y4bRtk15lGi8mLwcUb+TYPHUVCDij+vuE5zCh6RkVb9vQixs3ePfQnzSNLdxB1HCogFmu
XRMyh/6DgbjOTJE3TZOtcrdZ1NN8lVvL9Y+vnzo8cE+97eofYNqvCbvFgPO7cDSkz7Rjtu2rdl7Y
vSeHwe69XMNJbM97XX8RhxVbXXReHmJP7XM35ffO8xW4tDXSMyMZm+zJBBN2Qp0i5d6mkfQqc3Cb
IFUglOFOmQcngjR6Uu+uXdLRHtSGWeXLKt/mFIhSTZwyjpHydupZ3+Nn2qywQ5FoTEMcMfzW4pxW
yxmYz0TGMVxvvj7rAzBnKfyZizWJFgFSlX0NcdF5QypaMHNlg1WmBB6VBDCCRTcVppVk5IbPXg8X
M2z2Vx6TzXAgvr0n/mA4NqRXWMnKktzqaymMXNJ7W05OcS5AlIzjAa+glLK+uGWhDRSRGULPC7fz
RIeyjd+bLRmsOojPPTSsrmhv98bSglVaTqf+Q0Isyw04A9eVO6NYPHioE+pPk2kmdKgb938y2Sw+
453I0OEDRsZmXdf47FtK8HrH6X/JRRoEoIRFY3BBJzgvfFK2q8hkWnxqBcottJ6P1XSNb25vVZfw
jOFQGJTUbgF1lTxpNUHfU2Eki/oUeCbQQCErR6o3im6n+bQOmr+Cx2SvmruhGxWElYC/cMvx5xu0
jgo3fT3wu/fy3mF+UBiFOghT/Kz5JdI0xxpPvD/vdunV8Fp/fl4nX6mgTonsqnBHzG0d6ymWFld9
G+IXmaXgymB8+iUvcY3mNtJwIJZAugte5lmJ9yiegG5Vs93T4DJcpaw0GtIojbGKztSja/1xNQ/B
xNqtMQ495pZk4sKspOPV2AdY82tcrz+vrNNKaGEehlObZozZ5KF0G3jtVZiV6idYiCZHgmFtrdtQ
zBZ8jaoOdqY1pC6VymklGuYOkTbdxkqURLFGIMocNoaIU6a1JLLGu89LjjdGGYbBabxeW6O8OF5k
cVMXopUmbZnzdMTgwoYc/SPlrVxg2rSi0koj/1f/KbmaZu0Qqc9R+/wSzNWSlwn+0OvnbE+QaOdf
W7csiv+NZUu4VSXnq/v8Ia5RlbwZv1draxJ6eqkz6+Z9DZACPthaFpiyxPKUCACUHNRoaMQtFbuk
U7cerv1layExkgwMkRu5E4BK7gXiMjqLPfJ/Tk1OE5PBE6aXMqfFdN7vlyYjZWqd9Dgt5e/dgXLH
QFWqlpSynnJPd5quYM2QoBpQ0EshRYsL8VMM058PuZaU9+1u47mcoxacAhOKVWfb7X1MGZUG/aZG
QzORZxDOCFNldVPvreNa00or+6GeGx6yIHRpCnB7Bj30FiF8EnV1bkpc/a/xbExU8qAYPB1eNeCS
u1jmE2Ilu1HCYv4KH76vHLOadVcV7bVrfTjfCdZNraP91fYkay1AaingWABa4aJuPcOAy7bFTEJI
nsxlahWi+SeortOlKspcIckvLgTXPJjCmgvSgbGa8onAlAy7AqhQoqptRXnSLNLZLjQWHYl5gO5r
W0aQbbXnq7mSvLyu0RhAX3pK+Km9YVkas7ysqRh3J6r2p6yPassB5MFen5a7UJ/OGELUjYvPuZEG
apNYxDhR6SxLQIo92QodYm3AFZCXeu947McCiUwq/7rwMRYJZgZ047VyPWsRgGHUjnwuXQ9NkK2d
fH7gwmr9DTLPjalShM3U9N5NtCTfclB6xaxyuOyFwdQXlEb2AbMzHhQpku3b7haZmqdPaRdPaBFs
TDUZ1saVkEMYeeAJMsOxpnYYTWDc66YxPM8jldJjqZQLAbQfqhzInAvwbJ5LmxXZuwAQb9Xtk0Yk
7/HQ3g9Omd3ShnIlPhr6hvE+8ZO8bM+KkSXIz/194VU+0RoAVR63OeRTe9wPXep1uu9eGqg04Fy5
PJLZ33Rv7HR69zm05DYxCfe97qXNJHBqGJ08rCZK9PUQlgLTK43cjxbLP05PcrnRcKedE47XIr5n
KDd8RvCvGHacYryPV5liPlgqwCEWrKiAvqq7zW5UFP1xW+eqBv4ijqDVXlUv+Q1bd7Lk/SomvxZ1
W/my63XfJk/q6vQWQ5gxO9a7QltyyzmbLZ41UOWxJDr4BfdKc9QDT2I+1LRsYa7K1u2N09SEC6kW
GDqRzVNtby46YcqQ3F2tdSKytu0h+i6sq+JhxPDOAA2CD6doJp8jNvIUmJLGOggD3sirrkI9iGTv
sZwwmcyyt4wNIt55AOTKw+4jj2SYPqqy27qJqXlCDN7EM5SA04AnmT+btPqWXl8ab0y9HXm+IFSx
zyOobCQLmUh78FKFvqc1LpV5VFbVTI8AOWlRvr6Ju8JuJigSwW21WUbUFEKAqbV3aVmc/C6e/OcC
l+PoTmmxbq/LM6ZK353DpUfdjjf+0AEBCFOj3uyl4rcuattg6rcc6pniwGhX3T6RfI3wkcaHfi49
ffHpu2j954+MH6hW2VHRI2Hp2hQVXJDW8GUwHgkaI+Gy/AjcZSepwWHDfN1hgDzmgR3ZHK0wcucZ
h8PaBitXyAzZSL9UALyTIQoSgFb/xOnuH8HwcFz19CgVj+ZUCwIo6S3wQvPdFcEXTpKka1cH/qZn
i4Q7LtEo4hzwTnw6fzTJITIB8rlabMxx5+IutfiooDB2QoHqfp1L2I6/hQceaO6hqaS1PMhE3XFk
N3EM9d7zo7oQ55pfyU74FUfJQqZZ+WVYaOFL2EaNvDJ5xkEXgX2Wx60WgiaY/tZqf0qi2XIk2eSV
80TQUobWd+F1l88C/nsGxPBmqvPKAX8GuG4AUjgCXND3TwF9+xo4B8ZGeAW0K8MjpmcagPHsNpsX
DqrBGjAsI5qTOjAP6GA/JUXORTBoYbFnNvoTWxnsiI70WJ6zVWFAQ1c/wdg3zu0N3OC1lyaEgna2
skOHDbHeDLWBP8tXk9AWNZKzvRM4EwNMBqmFlyrgw8BCoissYU2mrJgpdL6P+AJ9ErwWUNjCJOMF
e24FbzwaHcf2G+rOlse1SX9ha3pEBgsPcx6UP0FiA3UHKtfjyYPpnpBWbSXC0I9AKHA4tqo2ygj+
ylWFuR/Tx2RADXDqGIGMKFrxhkJoBk1FBGbimFF3SufmGVW2Rq1ybxE0K/NxZb0Pty8uxsFqYZqL
rrU3FJVxionCPkjK5iV5o1p7lzqTyft7REjO59t8OBz1daswZ5xlNPKMSozehYZwVBx5lKEETfeu
xEGb7KzvNlTMM3H464EnsAzWmCg2D5LBStj+c2IJRoUYUVab/g3yLyhrX76w4K3k+xwDoRBufwlS
2WWl2r3BFhgAo5jGVexaNXD1mqwAUij+x2rfpurwT4k8FQY3O2gMlpQniQClnZjy8fm/bXRRHznC
zSAjKnqNfh6t369pHI95ZRgDe1a3mVD7qgzjJR5tObu01qVNaB8IVSSMeFNzBP9FfCe4cbIL7apR
xtgoVkdlFVbNQaczBbPTrqDVhaj4uqooGzkZpEphDerOdwQo2rESp7SeRIGbqIx0d4szqMRnbjqG
LnApg/pJOV72zmXOgKBrYWiQt99rC20kqr0oiuSlka7MjqOMliNpHmK9NqJxKHVnMuAa4xVyMF26
Te0mgzwnMEiMeJ5idMzNP3poqdVpS5WBpOhps5mPQ0w2wLPvabojQ2mO0BxTtAUmONo1TMvZ2ot/
lFsVuQSlRTtbox1C0s06VzBd+2wJj7zGlpnQdTT1zm1scbMZpk+YZdTDrlkRus4Fa1Lh/QUnkdF+
Z0qOJbctObzFVbAD6BhnDvz9e6cNg35GTuiVY7iRW1m2341TaSamip9o2xqOtX1hcU3j8uJt7Ocn
4lyyN/qXM0F3D4wjLPSATAmkEPmVCx9pXwH6yIGV/xd1yV9BR/agseedO+fJ9iMgFeB2QnJ5usl1
qLcfBwFyVghWxzDBttrS2uvXSZ2nycv97txIm/Ip8eEhjR0NTzi7sYDnaBZFp53ugfkVSiZ+2zVF
kx2HQpMMsJ7sacqyiMBK6U6Qvc3rVTnS5K34Syky+z6+YdHdTAOjlMCc3P5B9YLQvOkZyKDHNYCR
c9Q0Kg3c3ir0sijIc25oCkJH8U2I3cVTiNeuwDjYVKiGzuV2xSiFkkPjmJ9nKyqhcbarQmxRvtdA
9JIFn9fub6XWNJ62ZPzIiv2erlVyMLgQOz5YFX0k8hVganYpcv32tlDk6lJpwTx5H3SU7BDNdaYy
OuTcAK2WffTbfD8NuFtEdWJlytg3CqVJgFe1zkrh9SEYn9clfxeo/ZBnf/7kIECENvC4Ot7H0WGW
3Nx2zmxkEPSW0DT6qpse2wMIZUjvrktobibiynl+MtxDHiKnzvjlhEZ0C71EcGeR7IHjWg+yXvqx
lhSIXE0sNVwUlsliKt35iD/IZbdraAQoBCQvh0rNrgcV2Kxy6f1WYARI2jv49aPToeZaCdvwTUg4
1aivN0vzEetNg5HKKcyai3oEEbhyNXHxAf/RgFbLAELaOobapcOg/19psBWqcTH2HHECPtWazo7l
4BHNR2keRyvi+iJskWxBx/ntM4tEJulXT2yZYkfaHfakk/7JRDfjeRQ3ucnEk+9Re2YVyd0EZuUf
tctod20QRuok3yY1pGugcB/9dD8+87HcWfn1VtN7t4xbRKIhjp9Uw7XHS26Q+MBCa/OgEhT8qtik
XfQavjcVrekVK/q7pHHMrMR6NFNV6aSTuyNUP3xBsbU1KLPCwEg2VDJepjay2wOKUdmTra8/8ZAa
NKp9xzWPqkmnGv5xd7SCeUf5haitC1Ey/Hlp4wPqsGqORs2Zj1v6RAgH3F9Iu8ct+pxkYY5UosKw
g6ACk6Y9klIyFv3eZlZKQ1sXQaXlGBWhdaXu35QaTkWfK12Zvs3+T08DCYNs5YR+tALmbZ4tc99s
WAOIlMDw/mSuFjJ8qBScZNfCg41OGdRJtFXseEeKv/4c7PQQ1YyXYkEtMMc070xfsjwfJ1mLMq2F
VR7ZET/EcJciwptoZ3KoEkyi/oXQxJYCEBdf5bXkzwUIquD7NvF47VP3OM4H5ZLZcgXgTnh2uLDL
tazqY9JMdFW3v4Z+I6tR6VA4lFojGSrMGXwEanM9HNh3pVzEVqTsYtwU3t1gRvnjOh1n9FTt0M4D
P5RiIp7Dg7zEihEil4vNJi1kastil1qN2u5rSFcVcCS5JtANtzYNSrK8JAnszClGUdLW1XgCqKoB
z7AMl/83fBJhmv0KvQgByYJTnvO7UyT0LLaB7UAUDWD8/olLLH990lHUYOtA/tHMPoqu3I8uaaGe
jQMxu7vdOtMDrx/1PTP1dsZJ8gXWdWTApqw6fGdPn17HuUqvgUd4zWYxqZadb8qVzwny5KVsQLe9
ksTwUdl/DNH3xhwpbV/Fo9WFt9C+ztBX6rQzHUL1p5+0HmesyRdKXVyoKYLjJX4P9BKBqgO7PSai
kRRTLuIcV/HXEFx+jkTfgaXlLhHb8r1KpDwk7S8KCc3FhKu+cNNWcluEzEaKTxKf6kOUXm/EM31L
AU856gSwVz5EWoXJ6RggUMWfsHJwGCORsZNjtszpNS6T91oDqBmE0CuY67mHsG4L9h3gQMnlxNgs
cndeOhLdq6NeOr9Ydd0q4H7agVhObuJzJQC407Tsh5WexIjLRtYJPHUwaUooJePFHGXSZfRXT0/Z
0iECDVarp41tswhpfumSKwl537AEl8kiuDwGRLG288DUCGQY1zgIZj9W1ArAPAg/LJbk5wABFXmg
Kmfd/D0V3pBQmLDsfdWkXrPnH0MGs2WxNpZpaP0lXMEOpVQqQt/G1tAj0Crr8ValJKxYgGRjMinf
4a6FaeoWY39Vaoec85f4g4ho3U4ZVJhILIwDRsoPXJN75wpINUHd+fwaimcKGus87+b7+hvEVfDZ
h9L6AqZjTorPHjPGMHu48g0itKdpzROOq+DEbxcPyQe38VtYONUmVjYFGD9dwh8UpqQgq4d8HldX
/L6C9QZe5dABSD9BckvhhHiSWN3KoaKngqrGgblwa8RkuVSn3OipTlei8Oj0CftWGZWREJirKA5x
Qi9kkhYQL6UYhRgVv4L4LyATQv1l8pw1uoPHvJJ68IoApk8BUfOvEk50nTj8k4mdQWIb1EwtPXN6
GX4IoqWcpUjxhfFGXnKWUuQuzVR0FeTbdaJtB2udstVPUOXjCdRpXndyaK+XR368AauZvTy/l2PY
xknOgsXoBawa50HvfSLmAUFkE6fdT2fNoDZMdWgXrcsUsnA0X0t3c9gJJdQlNmWal9/mw2Rm2o0G
Ds/Tav9PC6ttr2alf3gr7mv7XdBbScGJiL4RPDgDDCrwVLpnXlbQdMv5Or5grBQB5R0mlJqnOCAL
G54dq1EzJhpj4hv//ffaWdyiiamgjTVTcgDW108FbYU5sDjQ79y0qUgV183oP6H+C2rXYOdreFDE
SycLGzy0YLwymx/ZlDs65RiwY3E6gBxQ7g+0WQHWQxvTFHf1JBlZNvbbESJa9/LhUVTF7FTUdiGh
s923qIM40VtEZNtcffDTg0q9PZgNLbIucOn316zRxPwG8HdcbXpetjBNTR5YXooWWI/OBZfXhpC3
6B6fXHD91rge8kSv7sjHNP/2/NMYizII0voM7vUP60UgnH5K9eW5wRbllfccPUSMkuYHvRraSbw0
s2AES05gKOVZ4AsG3FxUoZ2Midge0NoCmWiSeW/wc/fVnHzfAcwb8YeT5GaKPDRJF3JTOcAk28eX
9Zzzn5xz13IMpEBvFllu85kZ6/fHg4Xqsi3/Ou3ezREkGsEhw1CBf+Ho/FSQHIHpWmHO3yE8b3A+
yEv3RGt4IQmd5XoEVklRuXUBZNMmB6uWvDPdivskaFzlCTJAm6riNzlJrC0IyzhksGjg+w9zvWdh
p/93zTj7iGOx5c+n4mzhY0JvQ47OMiZS9quI4ZALbuJsVXC09filLavpNLQVBVPT6B5mQnAw3bRD
IfPbcFEHtEgkEm/hlugJF4+x2t9ohhJ34SntFJx83ogwqj+j5rxVHNBoBiLFSfXezEC+RNnodPQl
Ry9odorsLeJM+7eJ9KblqSeE0aEpK88Xm6v2doAeUgH4sBXzyXr/DE6KBSaLbUzF8D7SsPr2fmmH
TDKvhfQ52AAugEEhUuvHjZfO7L5Ku6rlsFnArPd/zjYWhU1me8pCxLQnGUDYhy7GC89mCDkanN5R
slCXrVUIVKlWrS0Mm2W+XlcIKdtmuRwtrG1HRAwbLyeRU4I703IWhzkYX7iGJBbE96Fkpx64TUUy
AtSAdzTyZh91h52EvXKWqktwEa/cKdJjPIyTYumaqZotpjazWLUAovVTYhg7Sa93ZDKlAHPJiW0e
xiZaFQ1EtUSgYwxHDzQz70qe+gh7boqS+SlAx/TO/nT0uW5+XWA3tKVjy6XAvb+3D4xuhl2cov+Q
msMkioSD55oJb+BqvowwGjLX7PBNP7Xiw2LKjLWnuFdt0NK7UB0b0sxIYR77Zx3DTUCWwz4kjp/9
8HLxYwqG90KhMue/k/9V283zY8gwj7RjIEGpu3pgZM47qn7gwbRb4p3qist1bl3WYmc3wikI+ESu
xa2gd8+7Nlaunp/LmOoFbs5K+Qe4Duc/1nn6GWZ2RTR2B1JLHnYR1g3OXBThB5W1fj3pYYMc5I0f
vd5xgrDVtmXH63Qft0idHpzlu2HolZm3FswiMIR8tpLUbZrn6bquP//r1RhuTIH2dFwp1zu8W681
RgSlr7M4Tn6PQxn1UB8gEMqpOY0PniwFJC0POFA2JTAeXeaxUKYUqSjxMQRCynMty2z4w+m355Ka
alBeTTf+CQXn9wc9pO0WM4aovLLulyrZj7vwLUSQFdilmwQXljkD5mQE/MlqiTPcW506SxXyjkSk
QAL3oEE2vDWP5VWaCxjMutLthg3EobJviLTC8ugxArq9jE0aSgrurp0bGt/Nu+TbU6xYFFBcheHj
hLKjEewpdBXkqkX17kxljzWDjBf9hZL5gyKyJDuXCvCPAfOTgBnIHW+1zrlKhl9JAjb5W6Y4Avum
ex0ON9u4lbExi98V1YsuNuXkNg2YvuBc12g/vRDl2YELm0Gfft35YeCCyTNenMtdNjiPNuXq5hD+
NIVkYAlzsaYRg2dB0MTSLM2Oj/wek2ec5WOltKPhPI8fBogLpDuSKD7GAZLw2P2t2rR+yVz4iNdk
8H1qTpO4OrjK0DaX0Tt2/aG7dAfsYVDwrD7yrjdjexBwaqJagVS79ia8dwhxHdH0c2NEhayfua0Z
H7BDkhvxnumsHZK+RAqCU9d82Mir5YHwgE6arMGSn5L7sIMVU8q9Pv+liPg8RgAeiLrK7gJVQ4G7
NE4HAjyW5Y1RR0T6Uqi9Af77Kxmzc13QVXqUyAAb9w5oak8Ry8OnjQV6D9gBM/RGwOtZu+pA9cKf
l3nG81/0f3zyIv+bxpr/eMGZEU1b3tERoYfexC/IM/8AfT/Omu99wSdD0DwG5x8T17OE9+IUKP7o
XFvG309ulDM/qwcu2QdJyuf/kwhm1oEmpvyvRK2tHquYs8Lkx4yoU5AkyMzL60a6tppOUhXhaRNQ
DWcU27GZ6xZQnhXM3dgKxRREhjIcfrVO3LvqBwHnRB4PZh2+Qz0YPE5jjA33c6tDhGefLDNDRX2n
+tilm43RPnw4Hl50HpeKZw4ymhoF1OWMbqm9sIkG8gErBYnOqSTXengt9jjYoArleUYzmHeCM/re
q0kt0OYtRLpwMlY/fdSihp94dVOQ043i7/I3wJYIcOrGZFXVsNxHdnPekbMcvABOg/BxE9b+Q4sX
zLSHBlVRFFJvLsXhFNESlodJ2XeDTUXbKNmzjUKnvVHlp3KFvoOu+EAqInRcsqvXthPq2obmbJ0T
u0tA0zvPlX+NwjrjosFbn3IbcjujImQSXFQX0psKH5O8ZvQgv2wcBkFDCqyJJdcmRLKNvdz+FTbW
3PV4WgfnT2enokG6oUvzxMhVUChoPA2z2jvGZSyefDYn690VvI/90eaOvnvPKegVGyi4KRfZ7WdM
Rfu6nJGt6JQtdqi54QF1pdYUKBaI2T5+kudwT8cYRqkAy8sM3ATd2A14L4L095/xb4Z/snzco1C6
t6eYGPvqx/SWvSkNr1kuRoOfKS/s6tNw3XXH4pP7aXAkxe86+CzmAuWsEhEnuzIS3S6NSrolCSPL
tGIdvxjUj8MFs9BnX2Q3Wa/taI5X+GMpWPtP4FtPiUeiLcLydTaov9eyDLUPp0tvK6JLUFmBNYmc
PyH0g8WvI4HVhU3H8z46vWTLtsktRBCFHH1l6uEzQp2tMTNM+cuR7KmjX0M9vW0UI6/iw32I81x3
MHk1reKSpTM4vjB8TCIgx+9EyCFir7cxucOal4yu0fK0RPoj0/T8xI/xa2OgeudmMasPgVizgtr0
yuPxul8r6mG+ECuFtGX8kaA4a/R+KtR82V2izprucyZTHANo74n9NRXhsj8KdU+4EyqG0Z0k57RF
Yh0koHM6jS2Oq8lsI+DR6390DTaVClsPTpSL1QLfSvumIosYCpfgzXZ7wef75HgTKhQSGqvT1gQC
k/zuMiBgRI+T1QsaSOiXB6b0lWbY8heJpCdkwjRMm63jxBrBt+LtakaFBoAoCe6c/nrxaDJ1FtPQ
1oPGzT+U6Uepgp9qOZ1hNhsCtq6kO0/40Rzh63Rxcl2okpLLi0jev1930PZrZndSe/yA/EMeN39f
mPvMIGDhfwfIxD9xbhL5VMTo7CSjB45avIyfaC/55+MjWHyJZJj2AJhErTUDQV+m6cRhAHPILYr/
r+zUKynHgnkSanF5CPCkDUXgZCkP9jgv/bk8WJTw/2FyAARgr8/SiM7ufDzRSNDTEbztAAHDRCyD
zYlvUowc6HgNODycqgWf2ws82uHF60W9k6cXr20fV0U7KjGgpdRtV2lWHvftO1Hp0R+U/pHicBA2
hZrW1n2+bvmF+edRKBvikC7OxdRtP5ygimDjT2tfzUU1x4Z00ErrS80ajyf/kIy4MTKIKqVKiaqI
89hTJUUIeF8+sgzg3biAMYBNutLC9PhjnUTYss9XVuOA7iT6jho564ik0RYrhDVcFdNpXLMI66EI
zC07Xzwjs9HcCK5O1rxy0FeNpc71Ah6Uxz7iFw2mwC5M9HVDsdEFl8UFji9lmF4WfCSVocaVcYAN
rZmvG5STzWLj27srNIQd0vBaxO5WJY3tnhb3eBBt5yvmzECT0jZLoJA+9ROzw89bac1+L4F2CV7U
RdhH/Lbx2unA0JXzBRH6GUJH1PyTfv8NwmTNcK2c1ZDPlpBpPceJQyydTdpJo37sSgx6l4a581WA
Ml2YernGnm2/VnmZay/khfvZ5J9MwEm5nZsU5BEerZAcVhO11T4upZJhUbOWwOdqTsRX3atKlOgI
7eKLGSA3/uBV/Pamuh47QIwkeG514kurNR2O4AeL9NcT2TCliQMMVpWZxJ+d9pC0q7EtKtsU12ZJ
AU/MHXZzCpXT4EGJ7512PtOnrICS9ISPeDlALDCyhtvDNpmJuHR1VO+Mef2NB07SgzuYDu2UAwEk
hxy3zaaYluy86zct8o2GjmAxUwCiXlrboyFvWmjPIcSLjAI7Epcw6L+dC4d8tdY4v0t0Ld1Dqa9I
ryuxMaQXdyzBf5Q0jBUPsyTyvbrzLjRjjzoBilW+/s64sNqD0mHFJ/whtoozb/o2/wF6VN4P+vmB
jlIE631tSGRALQHQh+JQinnymDx3qORWwC3L19mnvVB93d/3PYt2zYQRAEEPE+cUUtL+WMZjLl9f
HVYX8IoDIBSREVW+s6ViLYFUOzXbfdk41bp9Dxq4ZJ0oTfQgSAr++lz5b9UZLmM/lEAzIhuszMI0
nJ2DVjKIw9yENFaxOxrWY7/SWdYJL6SxFEUMfescK3uniL3qeDFxN1ltg4bEmJk95P9Jyfl2HApT
1Csnx+hcOWQuQYTEC70PRR/O4d+kH5UGOLKw8ii/aHUO0Dt4InOeSVfpVxdtpRzeeeTNklTTE5Nk
4LBeOCJmgrxFieL7dMBPhxa+dys1uRHRB5GYgBQ2LhC4yBd7VKUKUvS0Okwy42MkIdParOGSC1eq
D8QEtqxOdnmJW5WNTY+MUJpJaBERD5aFSalSPwJ+A6vuhVjoaNykVizTVRCTh/IXHLAGM6/5KqjF
OlTPrkNq94VzjIoFtH4g5Hm3fb6sDUDSWkGRTAEIC/FafHEFeB9MlftrIUfrXYlKwJGSzK3LGud0
9bOF7bAJGf8wJlbGX/dnPtyK3py+jTcGhISs3c/dKOL4vYRj2lIDif8OQ8SslMmYfkORv92s2DqU
Pj80C5NOKMn+D2+XvV3qC0PtckC4hRxSO8Gc9UAnGYKxQNMoOnuCGesBuAIGShKHucPMCMSzrTQb
hbr+CHvnXZe+pVdnJSNdwSST0T4shFTzYC4NamK606gM8gWWZ88Bgvcadau7nkpSfMwj1yxNQ9yE
Jdijj3nuvV/RGlXffcNhN73llc8zVnriu6BqQQeKURlDFsq3Qi+Gss9yPWBrFih84tF9fbjPKgMl
1Vw1YH1MAGyamt16abMo1EhdbqpNDbiDLWS+A0CdHicih8YJzQzcLElSJycCfjdiXucqZT2ywVRb
dPXvrbiQ2VwAPVsklLHBl0nVojmABNGagypP/iXRiDd72TMbYG8q/QxswQMEZKdJch/zeBDSWAs/
N1xAfGwSYJtmKpXPga3yGs88VQwCGPSYDVJvrI9AzvRkh5QvbrkD2gnwLhvV6/jRrlXawE61ucnu
wym/+KP/k4sz0LV1c0yYtu9MIyDviCE/L98KUXXBKmdgBJkGjOnPedBZsTpsV/mUNhT4RZayjtmt
qmIul1qE9Gr3hZg02GCUfeFYU4NLgsi4X+6uCbovOqvMMC8U0uMXk0DwI1ITOPdOWwhi2Hh6hqEV
YrwzDWdXpnVVmjCfS3DzJo0G1cYJYPO5LK+CpBtTUi5Wtxzd5u08ib5Jq6QebLDq9qmnXDWnYcsX
Dr/pLeN0H63BGpxoZW0kvpPAP/b6uKR4jdaQCfA5eDjCbWvQHcJdj9T6PMYBsIf36xQcQtjXCm4D
i5bsmqeKZl8Pb2Vtsb1Rq2v/xy3x8CQkfzbPkJnBL1C6FADIvvQzQqsP2TqEa3Bb0A0x2xDOkMG1
J3H/RhlXuz/P5BswoRhDUgIrdnpzKC7p8BY94nfW5d0bKEpiwDCbeAr2a+8MMrtiT9VyIHgTVFNw
VBarL62JbGBNOrVHuLHxNsQUuI2p05Tm7hbVatPVt3TSap+v5srLwyI/sul2cX+DJuJ/p18eR4rN
NQyKv7m5O9/T5fd8NLamF1lc+9kXpd5tiyN/MBLk0cpjHdG1j8C2uW5UYmEw3+n1KjYzu3rVj9NI
g9asc9j/CzUSxSjNGoViJezhxojztS+U6xOLFchN+Bv5lLY/TsFydSh96MR6U5C4d0mDFoR4U6wy
fIbDHIdFRvDypzzR4Mqo5Ke3ZVkpIZAO6KutDO8647k6ujQgCFRo5pCKFy6v+LohHinZxsXI1rzM
9CwPfbbk7PyV/gIWAwVIJIVph8UMQncumk/Dv0mPeinmEpYyagI+evOTDPau+MZyGbnuvhkk6+49
7gXAxBGwUmUZeDzZQfbSGktqfAOrNQWcHNDSyjRDlb9SFZdnFnCAH3cWipGgSMtOrdejzyIQUsB/
1jGGtdO6GyAicPa5X0xJmOixiYp76O/FQFvS9+x84NOSUXmT2Zp2KkGX2tD/RHq40E5rCQIibjKN
rcClQK1U7YRMgWRRodSOv/WWXrczBpKXRQj3v+qyOTkWq5lG3YggBuVkLcF8JEiddx6P2bitBxqi
tsRA6EIQf2kGYc2BiWioOXnAnTi3Y03A6R0rCt3PzQCZSrpbcM+nH2F1RRqdRVVs9PX0DjKHxuTG
jmA+67WhAUaaSy4siMbA6fUrEhlRmEuIjdR++OMWzNWyllYrap5P2L+pSIMl9umRTifm50Ca4Hed
6j5k9NGEnQiPywHM4hUtucLng0H0uS3z9Qh9ZZqta2V52vKghMMo/ZKCpVLJ+XIXPIXAYIRNO9Ga
drt7BtCopfttz0R/gV5AJFl4qtz0njwjaCEpizKKnTJFm6apGsGyMzeMAM5wYUz24qTzR2ROOZFE
/6GsJ2rdSSWK8zzndOLTkoiEn69+kOWoXEiOMj2R6FmDG55ems6bd7yhgUywNya4BzWpFtTSBFgB
RlKGjrKte1Po68/oOlLjxLflc2ZF7LgiQ51w7H7eAuvAmABYFXSjynLkbNEk7Z0TAirylECD3uXK
P90UVbov3bXl2VzG2y1lKFC2Mg3JXoBlxWW6Q46b1DXcPQ4S69GJHhCP6Qw8iQ6ne3rUgza1hrhj
/BC1eOhEuq6A5DCmKTPaCF7k55vV6Ch2Vlg+6L/CeUJdUBGMBMF4fFPMseOiblgkFtylcK1fk8rb
zTxBl+z2c9a8qjKueaxE34zgx1eNSOfdRA5VSzo4W7NLrFmWdd66gtWsQFxpv0JDJphd6t7Pf9V6
2EWrjN/MCXDVf2taS7NsVNeMb3owSXx44nTGLHlqqbqzb98VmEgizRRcmYixQFNdBuQkPwTmCf66
tlqffHxkFdg8xmrPb/gts9s8OAMKLOPQAdGlXiFQrBa3jSB1gYjDViD/WiXyeXUMKHKcjzworHOy
hQ3uOZSBa073w9cZzCzb3ERg4780muqdggu2EZ9LJg/dW0Mu0wsAXRtGzVxUs0hUZ/A3BsDUB+Vr
8gTgxjlJfudeB5anadrVbDExUf4C7u0BNI/wYZvrGwf706NkXr3MPLOk4py8Fd8kzKYNcQ82KFKh
mHA/IOepngrVTpFbw4qgBM7qKiZRhbsXf2tYkli9KHFYhUiKmqkKlDfUdVWRhaoZx35lTozLvoXU
G/yx5DrQm2bC6kO/RF1SEy5NcRfq1JPNera5ScT1gRM+CLvDRS70F7oUYbAcU5B2svFcRBosastq
Wkx5Hpn3TJeZYX6O3czxdgJuENr54OFvz5BLtTtR8z3hWTSMOsTbFOWd8QPfFqxXHxPl6MHnGY93
7pdZ3fg8hvgY49yS+ddeAfDPA+QNZhOqsUXoo9PvL6+KVIkoEHWgG4YaNcBrsY64/GXQzHOH5xQr
3/Mx/onSZWPCqbLcEjZsDt2pHDkluqzHj60tknjLKlvf83rQhJ7NRAEztTra8cNbONhSPA70wcue
rZMAERAeC4BSDaDpDklJ2BA76X4ClKzEth5GdXUUc9wRBHRS48Y/7HZT9gbey5y+X3F4i2fsblSx
TvOfOUfgKHyahMSHyMrhhoRS0HVdRl5KBIEluEwhr75M+lsJua7bex3HWgA9181RtfSaLvn6m140
ov4lEm3uhLjwShHydeK/XjQOVsCK+voFqgEG77pP2Pq/hY0ympIUCCNoTfGqfmDNKTZcNKmD7Wt3
OujnUwxaqgP1oJ0ZlV0VD0bYR2466ejjJg6iCT46KxIu6UF+w4ybOqZRRaaEpppxHOQU+0tTq0g+
W9AUVkoKpsNOtua+XRBYeVgtRTzH3N4rmeMd/jwvgGSp2SxN8DY5Q8u2yevs39A49g3BE3KIzx5/
ULlvkNlUnVPusutj2NiU0w8GSOnC1PBl33YnSt4CyGkCzD3KTROmkhSrPniIVqtql1zuOQ756E19
Bbag7rTFq8QahEK44+SmCCLJPB0YILt1H+d3nClmLIkKCTFZG9w/dAwOVVkGQZ3BlHVq2wi0GQqR
S9TD+hJVsTU8qbgfH0cqOHm7DCG43WrgLLQPn/kHKIY+Tv6RM3fM/+f0smRzTgWZZPKpbEYTXzH/
H2Ol1rUKsZaBDaPALjb3e2i8h/aY2/3pSu5Rry/PgxsEzG77x5bxotjhB4TMVmlBZkltN4eXN6eY
E0+/wGjJ6qIjB+2YFtpsoD15OF60lJBFTFLyEUtosXYWMyLGfWa1p4fNyUBCLcymab1/upzMDZe9
yWREowdOCGmrcyuE1SjaSp7EmBdScUvAyFFldDkki3xqSlDlIzs2AaROLLbecSartymX0fVuxlSV
qTE7YK4sTZbVfFD1RJsohYVgGh2YSVbQp8Q2Q4t+tpRZ4uLK4/k6dm9Fn/upM8UpeO6WUNouBMF0
zbfwb0efU/2OnhQ+JsvfgF9wA8lQ/iWxMdWWAeiB+qoABOjb5SC/5BEeHVOWDWfUP2+OYnRxR/Il
ZlPjrfnWM0hgMlQimJ/6UUHkTqdWEdWYs8m0AeqwqUDjMt2Dt9nVyOGCXXc7hVb1sVQ5Xrmwiud8
Sg2vqYrUOo/RqlQBgWf1dxquYhV9551VRjQ7sDK5Meb+3iPRBd36mUierKrcC/A1q2cciggbTTso
KAIwu9SIKzsm/YRGTTuiQZUXeO+yxuWigQaBykYGbz/VIZJkgZTyQeKFu8RzXNwnvfwj+8VFiSJm
K5wK+KMcA04jA+K1DB8cP6O0Avg/hAsxQzeXwz2E2L4n1bN9TOPb3TWrosREOPSUbWA1qhf4E0Ee
7iowbpemN0SaHBbYTKg7GjF1x6Oe9BdHK7d6bPgv2fjELlErTWEuTgToENsofy3HHbzWIfjVhUV4
inOpr36fIWV7CyBJ7ofvJbFyafDB4McMvRqKVELBNegPePdAwSHNqb4TWNLYSxWIngLzifkzjP6w
wPuYuH3smFW7j0/U3CPRARGZSs/nYN6Yn3DolA3yVV49A1XwRFlcvx9IP6fmqhxvlkSIfi3k5lTo
OsVsqb8ai0EFdKS+hlpYi3A9b0tNmN6Z82ig+RBoZtNaR0YPK5hQ4onMsrzg5a1V1hkACcZ2p66R
K4n6IZvRTIQMXOTJYzw9VqRtUTlndyt3g7Cqsq0d58bJ/Wji8lGFtYwcaihXtOSCYpGJN8Vgrj2f
MVJIja9JJPtrbGmevWslrfN0hhvXl3pn4V6rQzeTYii1/Q3WJ7nq9QOr96+eMsBZ9NJHYXr238Wv
tdvytKUv2/IL0+7D+7uwvCcFzDq6rTZsXSqZyGCAy7PHMJgoEFnh4RehiTQryJxIHe1K0LpNbG0l
sKyD0vkr+4YobMQ4CTdW3efiFtvsqn85in5+d60/EJx/xcd6DHDSPNGh0FY/Y7lsMRXGPqB1bF+/
vbk2TDYvaV5idQEZ7gpwv26DJHoNX73/6+Lv3hIdxfgyJk6rIm1uFYG2ECtPdRrw2TJRMsPAgzwP
ZgxhKu0ESNEcWo/RpbiaCX1r+D3EvW/rl88sNRSX1ZXd9Q0+pG18OVnxSL6pugwxhmheDWM92hzf
g+NA3wFJYjo81kXnCxkUI2A6lCZQsrXsE7T5RDIMR2X4zgSTI1yzGrbZ5oxK0Vce9Ql8FktPGoRZ
4q+PLcNiLeq+S2CXGqEjxI6pYpyoUgkANwCagvxLBbSbA4wr9WPf0y8BKBili6NlBV6NMz1JnM9f
eX5RhnWrgyHdtn3SzKVVgmqbCtuL76s9uUjs0QJ8MmCB1Si9/G4/flkKJQDmDg8uC8zFL7fgZY9S
cuUe+z5ZEfRYgvdLSLjJQ3GVuRxK0JVCPCC+opMIR937+JNk1hNO11Xy9ed3dqP1V/30w8lQ8G6o
mJsq4rotapbRZhuIDtggkeYEp169PbKkvWHx3Abrn/afw8W/KaCNk/Ks9jk/SQyc86oAHWN5X8+w
jDOWDKXoqLcND/RfhhB3uKz6kxs1deTVxEHjsfxAz5NGNO6rHUxV47O4e6Xr+UVjW3PjSFqMVjp9
rjwr0KY7jE4bBXuIxmn3UQWzs88/W24CV24Ionlfczm5QTYSop8KpEmJCpFikwpl7TGUHVYPj0mB
MsEb7nLxP5utDe2jEiWo0mTlW1+8/ROoQCammMMBpl7t7QCZFXag0rTcUQh5q9cimuKuZdOh6eSq
M2pZtcChAXpVnqztVH63Wdpqh/g61kUlOi5SQvtYROeaD5eB7jQgrfUeeQnkNIovZ0s+vf0glkHh
bhEhULg/2Xh+n4OnWp6AUTO0Kpf1DJMpvQ7CW1jAxnRM6Ma6Eqkpmkr/ShWsJJG333s5C7rqJ3Qn
ltnM7Z7Lf0QDuNK2Sfae9SO3oy9rohRRfhsya1WXCnN4QJsvarnJnDYAOkml53HJZ1C/x9UO9ocF
7AI7IJOGx0xheOBdm4UxjLJLJ3gkKwH23Ksl+emRiZ8QQPiNooAWCSo3xeDkeNQp9dO8yu6MjGA4
prgX0OzjNH621lBr2bzlBNkUnJqy87HMMzzqsiO+zCaz5/h16D9Iscjz6CekY6DpRklW1N89s5dB
XGh4BVfhpWoJHgxbecgX9gdrlewtnijbxCrE9h6wybESQ51zz3E64FyULx5FgX0O9r/Wvc9q+MXb
IPamfDarq3m+2oJSCFP75tejUxK1exodtGiszDY1zTjrLY0xgmPbU00qSsdViCn+JvVPSAnyL9/N
tjvxMDnhe6UxNmt1KaIA5gB/sFQTT/4CCvuVNkMTGc1bIMtroKJCUZAKtu2eN1fpuei1EGy3Rp6N
GTzJNDSl/XeB0NRcT6XuTStVA6xi6q9dCqOpfohAS5EDKq8AehwxZqmJ2o/h9wBQXtJOqwYy8P5S
95fHcaVAn/VgwtM7HgAAvwo97TjZD9k4qNDbLcRHGMoRzGf9khR5+VVaY930yDJ2jqXMKA7vG65K
SWAzZX9x61sOn/cThl6oHAKFZSHbXy/Nb+KfvPS8GdIF+nM+GLXy/XhV9Wh66kKc9Xsav+g5GtCv
q9VQ7Fgh8mUvBnpyHCreJc/3Pk3yFyONrx19Ze536owr23sa54xQdzV1EoGiACYZb+dL76cvoqMb
IazhwNuohQ23NpiRcjQzIA96pQT9+filVvzLjIOa1QzwFKhoWht8x6Y/GkfeV4agEkdy1fN53rsC
lDeaOXOGm+pKPrDIi4eyzz0T03xd6u4iM6URkNwIxqTi4mbZTyU0tn7wr7JeHzOCVBqEljFNUWSY
42FtPDhIT6PQDlDZQOcOmU+HHGBrZPvTLzpr+GLs+N9gc8YhmOBoAMR9/GUPmnc9uwKj9jh2gwjt
1ZF+5pef+YVdsGG1w/6h668O4YzvFF2lhsrjefOEn/3XHt0oQAtNu/gJUkUjqoFakMk/vyI4y3Ny
j/Krrm+jcP1dCgiYfZz8z8G9JveC3XmzoNRgRGAoaFOEC7KxY4XvGZrsT66msQgvmk2X7SXtk7v1
PqJHLigS/TkOB/MyYKhUMCD89bY10I0TcukGtisxtcka4d8qECam68CB0cvcY9qlZfCBhcguSp5w
7kL1KP7j1PcZj9asXY/QNi3wPneJ3WjkglgRbCW7kGYLQioQ6xcBUxpUOto3CAc6vEzWVWcGUAun
a+/8aYpZZkKukNz78pjRoRdKougNKHoeBNfJmjjr1+MqSJfDmGKff8810jLM40eioAUxwNN5Jvvk
fvldgL/qSzfn9k//j7Ay1sxRzPXCKZFKzG1YxYcsvJ0uTdRGypzIHtkq+yM36FoM/qWUtcUKe2T1
UKeYF3qBXvJ30Z4vv0ZCr9VzQYHBdYxwZRkbsGDWCTFCxzBMmjpyyCTikCi0UnEE0R4AzQRdLBUF
B/H95xDbTkhcyWNcnOATi0dpdiGhRgTA9e8hyYdjBCpZhiqAAy8Wq/JD9xXuRCfNv4igElWca7Yx
JELvj1OyoWnqTz6eUoh2L3UkaFTWPKLjMobSG7NITixfTt8auCUwTKsAfQ0eZMSjmAD0zMzT9q4j
i0p1/bZs5HOTO0/sM9pPtqBaRHwR5apiDd6JQSoME96Skp4X8ESAjchqYe5UObFZBKUKWzDiP8kl
I92fozdXJDK2Lcwo26qefzIs8REz7Aa5RGtq3knbHOI6Mm8Zipq/7kIF1IWlrLy96LeHmP+q5WLa
F+ZG+yZvtDOYvze/La2855rd87rVwAI7lJDuWlFyUiivo9+8UqGknHBlKET6076zCLU/qbX/hd4L
oO4wZlyofpnj8HELipB0aFl/rOzan17B4e8PZOzvoZwTVLJouiq6AZ1rRV9q6ZVtbdBq7w7gt8P7
GwN/H0ZSxLfCW20Kk4+Y+IvR62CvJWxjY2TVpCwKy3zTK3SRDikB9IRuPsR+V/Q0SIzihJqVMjgh
/H6m8B6E1A/xgTaiV933dq9WNU36NME4FN6pFhGpNfoPl2uyHbzSXJNNN89YGeHQUz1OxOK0fSeM
+ipmpkPtNFMJ1OveEbIDIuW3l/LhZmDCDvALa0nbN35/Kda29MGa7he/7IFDlODb+4S9OD90W5T+
8mU19aFpVcHjJYKa+OsRlXkREv6QZzASc2yHlevgKY1C/5eN9Iw/Yfs7Tonw+8tCamvOp4vecqz8
OeT6NjYat5v9CDmWpYIXPxJ8VjpEaR592JK66jtEzT8tMQxi/fsJTODk2Jz7NqRa8Z2LopdQPHMB
aMXRBmXYKY3i9pcuOvTmFUJeHuxbnMEmp//A2QV75r71g7CtB1BUHBRSjgHFF1wASGkPYvTfUgn8
o7gIk/Ibl6sg3rGfKltBRtmLmgKjA85dAa9y2nG8Hcd49KSNTdKV3yJ/MqBLpJzXhF5AgH6/MHsm
X2iOwdNHI2PqEuqACiKNu6w3jyn+xq7ei+2FYu8M3Vm5qRCoERXP/cSwDTBsHO73KVQJOJMAgcEN
Not9fQg6+E0huvRUvMP8gCHZ+AGVrdQ2VRrC02NrvJCPDWh2ZubeDLcokSGuYuCj3JEZDd14OkRi
GbE/f3M6IRkVwyJnWk1NoqXLw6x4qos3IVgCs+gIH56zLN8zOsb+oq8YHrr0W4yBVxbzgdiZ5RV0
voac7hHr6QgHvMdxRoP6ZBLSsuaWc+as+nF0PAl4ozLi0+9Qo/g+BdMWKTUPia6OyLD2yzRZWv4B
u5W1xq7vmfHgOXC/n6FWVFHX0tvZ6bmp3tmqmaF5zVZzimUQctJ2pGFODubsdRrTmzgG7A3tuzyO
GYEGXrheQCWoL7HjUV3vuE+5dvSngHyIbZAx3HJ74qx1F/7hFlqqLZrpd6kz1tIf+P7SQn7HTY/8
qQfDnVXEMmkBdOmNNmo7hs6Alb4EQZgLI/qMAujMGADAREBrjGk3s8q8wwjMW06z1SS/eu6IYM0Z
DfixfGZ8l+pq6d0PjmWZnUtAKWS+6y1jlqAoX1JUMTlkr95WS58cERRq+qdiLvAj1dOt5JBj4944
kOXvarOpYYXCFgxB3y/f8Vx2eVeRizhm9QzGkaxe1bWB5TOPTWbvRUxtKczhkSChtf8ybjAd1xzi
J9UR3EL9f6DxYZ581lx8h21mcpRBVCrBeoVFVvqiYyDEVWPN3uKBxPu+6yQmCPS5Io67BJbo9KHC
aUFyUi0SGbyF8sO4N4kg2NwecxGavzX8cb2n0w40lpSMwgNr9f0qjGY4lEDgT7UAiJcoT66qHq1A
64BaTTJgoKRQke2YxEEimxW/bB4yKx0LEF9qxJemg7DfnZscX5m0nrrAz0KKvdoMmsRr02QFw4q0
hazoqYFj5nnSf6truOvr/jYGWxqykwTgJef/STDHPH6Ok6kO+gc3lv8hDhbVOghPmrx4GS5eFuyy
ZAtxTVCHn0JfNp8yXs6g4BqpZPeunz5Yab4kF9DlvxObgHdbTqW/Qu2OsNFZsTWhcIvNLfEPwHtc
TOu+5/lp8UBdRDJt6anwLSbC0BI5wS+Ck9kW2yCmehHR60dHXsvPNisdGS8dE9fRlZqLkr9rBw1s
8H6wweOnNc7tnQ9ZN3fxT+WE3oLJl1kGknYJkmS8MOJ7rDVMJCg58kvrfUqn9OPhMEBTJL0NINzG
eQQKTkADMS1pm9j0ODob5XiGV3AcOyM/GL0mydQlEnVbHkduUhKQN7TSC2JDKXT0Np1CKW0eYy5n
7PT7YQrTHksiO0KfGV8s3w0Yq6hP0kqSKv5TUPuaEgcOB/BWA4ECxV4AnqWWaXcUmi9riR7XJX1B
8cd8kOmOHXlct2UHkk5spCqBTKXiEtUzntvtsECmMMNRnDioNF9N7AoMk61f7pVZHCgvVgYBHfO6
wKPy9qSqbCWVVIkSjtOMK2MZI8Ah+zqUpJaMRwbcadd2se6sZaxTQbbpnWkMWuh0CfHHHzOy755/
fCHBQdC4RfiS5ES0oGPj46EKafZx3wsMCRvPt9+adOysagwKvwhL+v6hAKKGazM1Pl9vv7FgCGrG
aj9iX6dNomwLXKWiGHQ25SxC0Gklhud84i+BLqg4IsDTPlIomqkRw0E2hc9ux1S9M6BIG3/S2iaD
HnSHS+wrW4RBiUzIOiOLvLwT8VpDHDFi8CnerinjvmcKCewltv9xIWCRZ/4Ei/pcYPlbjb7oy+YZ
97z/0zksIfn/X6PS7uGdisxHP7IQyz1tLeHLmcgtchkswYe/7k6SgxjX075WmUYaFBKxhKAMsBmW
nA+PoZRieSmP8J2+W/p76bWxGSknlaRBhMOAxwTKY7q3rl9jAVSnHOiDKnjwAuZlsIcLEERT2KKQ
MkfbBVLpHCilYZa1XtbPWKpEm+/f3w/R2HHlaSm9+eFdCNIjbjK9ScyfVu20Lgx0OkKzU6eu786D
Hcy6Q9W8VxirL5fe5QSQYj3eZFlWuhLNHZ89A0IekRBLm7v3vqrPC0xwEkdHXn9fnNYwCYzmlDCM
e4x0IlJPs6dhcVGNzll7tHT2yNZ1Qn+wANE67yhW8nKVeTWYTKrmGIfelKGDsk8uGCUrgq5drBne
ARrbVpdLa8kL3PKhbpH1yB0zmpv3JhGo0s8H5hQyfhcJt7Wf1OTzeo5jZWgNS7C4DBzbMO/L3TOq
g7Jd+txjHxRMsLZsbnfIOqp65jKbWXHstTdKlxCG6URt9P1KiMUMKlNPnjdKmi1GaBLmy0Zknp09
JJT6gZi2c5ep7LaU+NJsTsun4w9yeqsUm+TCAStmd7Yz/LPOtDw1YOo/RoMvd71bx0QylUhfmh9b
plYP/sCBZ8qAAFl8i1Xq1E/BEPSWaA7w5qXcG8WM/kNIw32D2d8/87Dsa7z5VrtUcs4gJWDu0HjA
NDYzgqwS725Ko3t41L3hmOv1i/hQ9XpGpVlxGPNYFHuvIyxY2lXcGmD7/Cw3vxdf5Gw9TrplNmeF
wnRPXcDzh5Kfi6JaIrasCMr8MPsi+dXPppLNq2WC9ESW1AYhciLLLiiSkDRiHSno3amJL9AG0ck2
8teJUAhlTkbvyOK/4v6vxaNLPEgz8bquImeUyINNI4WQS8aZPppqpS9Q1ewHphBUGMtmpcIKYwLp
4nQUXRdRWK+ACHprnsTG7rsD5vOOCOPOpIFytmIwZ4cDZIQpRd4/wJHZpn6zIKH2/UvMOtl/7A5G
06cOwz+VWpFLCYVkfD89CnHGV/Na1SNPcW8E+U6mBApTsw3T2jT/7e2wpMs15Qy/sT+yWYAW9Hg4
9lg7T6SN2YPf9RmdWqSo1UkW4yhPpR+j46K439ntq9iht86rpYzQY518pnyJVhyPT1Lu8HjU3j9V
RWXg+s9yc7mn/DZLDEX/Tz5ck04H/3Yxydqlv1ijPH54/2LoDk8v8NtuZ3OhVo3rG/5+/CFZ2bi2
nKX78YynZEDYeCB26cbTrnxXO2qwXfV7+7HwRzyT9yVveHP5aJDOrFBoHMIexCKnnQpbupiRH2h9
1qQ7IfMXlMWpReLJqMNzv5dkp+o+d5QpyOjy1V//UAXqh6m283sAeEzmdRRvCd8vux41mu8xtC2e
b3RerJq+dOBt0Iar/0btnZBJL1DLM2C3gOkz73PqKxnYzfNzPGbCHbN7ikQ/sj2zI827j8A/HZ9F
xoqR6UeWwLWxcItVBl01GPe82sLY7znfYAroL4U1RFuZTja8BPAmuB5e9xVUEPwkIjJpdAi9pUVU
86k2XXCd5pDkjnMKdhkLh6B14dCWdBlqGXb7wJ5bk/cnu5Rvfs33/e33R+LmlrAX16ecNYUTDS+u
AnL0ZeWCbGSslRoUJUn5/sTNBeZaC+7DELM1SZbjs/LCq169Hq66KtYzU4owmLg5g73hfOorQ1a7
HiuK+21uHowz3C4Zl1EVPqTMPC81i4R8be3TfqLic/NQe1V3wjm9RyAXkdH7AW1hGeRoeKdCn9rr
64oFApMtQczVIqUxi8UH0t35OtZmNWK2c+dT9IMVOCEUtjbZv1OUZfh7kX6Y8clKEjBWn2HEzu62
TYchxyO/TDhTyKRv+xe918rCZapW1VuHrlVjeLcTvIslzrIj3/FU+Pcl0sEAWYyJLrE4XhoeV4ch
t7C6nEPzV91eVzyTVLruTpn/1168+M02NJwQdmBmLWylBKK3ON8WFYqYR+f1pPmYG+Jlpr5Ig1jZ
foXDnEDeHU8USwOwh3tmKJcj0RtKK+X0GCXb+CRca8sVVrRth5O2LwPFnQpyUDSZGaHc+AbZd8sf
FqVGpF3COQarMErBDlySJt7Qat0kbdJZirhy//atpKv1dee5iiVLQNw2OrgIh4fAGXQKaJUyC5Kn
Fq+u+LuEgLQtZ/5ra7UZ04hxPio3tKYvt2G+LjvAXDEMV2SDIvsrqZxC9/CuveU2nguzxIr25Mge
52T/ei0/rpS2NiClfeuuZ1x/Pp2+eKNokV2DJbEZ4V1DfZx5Ni+W48fQPopx9SgA7bFmj8UZ77UV
Q79yaFYlT2VM/gy+k09CfOEdEosRCQsnB17AJREK+OV4ky7C438vOQbJ2c+cRI3RYGmSDnoLDLsz
oLrFCKYxeW4FaSKuj5ug4Xyva+mpqkObnB/MkVIH7mVXmqlZ9N2UtX+XGrbNaOjHzOLhaTJL3JP9
XZjkBIYgjcwdK6v8bBV76kUaAqrLSZxoGujewJjWVJQFY8J1VrbymZPktqC8QTvGmefoTrMjirUs
keSoRJOwy/EOna+DsIdH9PjfVCFixtTeMF2vLr+/0mFXy2G4DwyB2z/qWqH5Fjl0cx+HIJt96Rn2
StawvyMWXSvNZUW19Ng4MLZTySg+QxbH2Vhz8KAg8bjMxbumEvl3SlH+ngM8g7RZ3IxsGCx4OgwH
zUmhAVaLoUX5M2filsXlEj3vRmqx3eTfFtAh1PKZV00UUjn8wniGEw7oOaWcVpXgZLrUlY+PJaZU
neYPHUbD0RZwlPQJc6SdSpggMXLGKEYPWwNME2Bp5ehW6ZTih8k6+Wp9APktmm49fovu8yk3WnKJ
auQ2cCPVzQonDpZG/Rc0yDnAVwm+Lv9ZuQiMdDJSU2KxO32JHOFKxt6sn8KYRlyNg8bsrar+KrKc
8UcYQpBVwgdAVrTry+j0031E0NkKBBN4KSI94aYVidOZ6NQr+tjn6FDHsJBAdECv50INBSG1TZDR
b1+8PlRduqVSZZVIDSA8FnO3Q5h22f6w4XyUxXFaJ1Q1dytfqInN5JDfdE2JmwpLklV8fdjZBzzQ
KEFh0yqo0bMvLW7sAJpB3i/Yw5BcqJBURN5OSOSZteMrWEgjEj1c8/LMGybDtwt9PnWaL+my6zOP
POTru9X3oMYul/sHF0yjdrkL9cZtfFVIz5KAW17NR+jDqtSKWjuTgTY0VSQaJpEw5gNzefuKrqAY
NsDOEo9YYLYZBpeCtdfRvypqsIMASEWgjqrZxOIM+do9jcJMDlFoIYSp+SF0RwTfYQLZQfOZkMhZ
F+EWVgvGNCTf00BS0CE+7a4RyzMVNUMZZ9sBvpE6RHDrDNiX/JwwCfTk0tSlCItgSaWU1oPxWdEX
wanfxwQ6YKsfPCIcMj2n54NLFYGCBvL3kzJaJsdTarH6mPx6L6Mxt0R0TrHVUO+RCvBAIicACy5P
+rbwTzY6rJWc2gDADWCs5LJfUAiMD4E8+Whi42N8V7V9libn6RcYH59KTqKggiZHnog1HG8N4A9d
PyM9QZJOJ+LaASNHX5X97S2oVRagix0M/UkT0Qvco/blRZd3oLgjNZ2VXMTVdxgOHl8fnTYPBD2K
efD7kmlPfJ2p7/Rx25wyXB9hyEUot1bWpqElZqQK+GQiMxIB5YvbS7ejKM0MtqJ8dsW2G71wSP/V
702GULm4SXAGbjY5tvizqr083fhF34h5O1oJnoilTkvt2h2Gj4W7i3CUnk838m9ij7weMfxu0z5h
W7ExTIQXluI5SVDSPCH0/yUPmdtzi1JuSTcvCvKJlgYO99Wu0XieBEYMJwnuFq3iHUTBhBaHA5RX
Wvg2iN5Jachrp7ALAG+LsNDfRMxiu207Ejxb34PdeHssMSHFsK+Fp3PyJZCMLblpp/PA8s1uoIN9
HtsfUi6VLKjM/XlobSfyQLG18y7O3crBXz7U96wxo0zahlzIxP8I5GXb/6tY/vOA9d/11USKBAs/
SvR9th6eXQ3zzrFxn409f8Uz/dDILt593A+CM2+YRk4mPK4rt3uI93DnnTt9xdD8cVpvUkK4FaD5
FknXy+yAK7lTywojadxis9dXBNQNlCwjxA/7dK61M5Z1WYsbkmW2aLRi4EFwN2dbQZOstNr4AC5m
d11yq2TENbHorHRIhOHgfSqsdu5al3HtSJqOCVGrmGDQF1cF54r/I1T25GY1zmT1k7Fa1oKL3bFc
ZU2/is3rgwp2EjxxTgGAKIXYAmFgk/uUq8/jnjVmi3uXbRobfgnhcNy2TjAO3bhZWORKaYtx14lb
2HgKFbj+/YSHlHw2vmox/NfbYD15dx0QjyPy3dUkaLPnSZPQhMVmptN5u3eIVWC/lvNcBtgx7Lnz
iqIaILx6Yf250Qu8PiEJq4XJks0Krv/sJetBcCNgPbIVuwwCo9cedPdkTDjZyS+JDVa2Tuj9E6qv
BvIUnKN6zQA9jsZ7NN8pa3zsaxwo/0ATf1vE9fu+HnK+U1s8Cy4IvPtRehPofjehKWq3GeQKUrK/
0DldLy6Xzd0G/PFBy9gQC8lthlnOacjli4fRACBV3d+JidUOY/zT4aFsgMk46oiRTg0vJg6wnCCO
W4vKm2yFBvpfk2ljJWOSC5EuPTx9BydvBmpcxAjY0soHNb0LEWxOgvl3+2fl7ZQw1CcnXxnvILAp
TlO0bQDKKBSjv+ri2bHcZQTOBsht5DndLFVqwhBvBAAGZhnoUldBlzcfoutapR6WygE9klylHnk4
i/yXV/3rzIZcAoVqz6Yh+rw+nrWkOkr4G/Wj1PSqCTgwyc8Pr83DtT4MvhXPiX+3lMDkP/sCEQJp
+hvZKyVF+Dy+plJJnPIvByx6PPKbxxzftpZVKEAQAGoU/5cyQv+j9yuq2kHuUhfh1jfpfCD7KzEh
aIiIZxsSPLudyO5rIhQb5N7yPOFdoAkVKhOQkqEblHggHq6b5Zz/e9uY9meqNGsQ9PG/WG2YLZ3z
9L9cTON+fMZ+WZOw60uVo/NSSicoSvQrcko/ZfbhGzQMCutzyb9/n9vasLYdsxcJ2BZKAONx00VP
PXMZdVWkKEJNEUzhdBG6yGphPBGTGzMl+uzAYexins5K/mwALDXsj/gtOMSRzxlg0eL1x/r6zteV
zmCyzMOXLZ9FhDaERUTk5AKY8PJCsdMPyQAySp91yrUYDQw3ts7R6WybqgdrwZkITP5qAEYK6lap
bZW2F5I1VqPSzaMGqPLp7/2pzqdeldiWPB8jw411Lkkzi64JupWFkjV0azSYTBUCZV5fH1LHAItc
L+DYRsBwN6eNe2UGh5wHG4mag8AdneEOR2ryfxJSAApfNZbEURxWaS93etXG0YBUqZohrbfNiYdA
f1bwlswLBvFCq3bOK/f8Dsmd/CeSyCBjSpRDw4mkK49ZhDBA+0fvozclUT4I7TvR7lQ33sPdtdlw
LEmMziMCj7TMXlPolECW1Snh5adgZLjTcZfM5bDT6iwpZC1e2Gw+d0MNOjYc18Xbi7mQ4Gs6c73k
ZJrM9hm2sy9k7Y9129ULNdLs7rzqHntCkNt20Vm0l7TDD9fgPZ7X7Rb495AEFLtPVX8isVEZ9ClA
tUNtosc5LcqMVo40hOdbSvkQd45WQmlf/kmbV24ZsIogdCEIZdwc4yoaddSmOoFwxfojlCtnwYSE
kpWdWF2BP2JKXCvAuYz61ihXT/UqwuiULZ497vnNC2c/ED8UN87CITveOdc85aIS7X3Rq6bwsAns
ZjP3vXTrPfcc8zL8sqEaEJv18ypgW7/G+yZDZ1ZFIUdElaXs9BX380gfSrwtdwfmFtHCaVTMGZN4
dIPMgwVc5FydXjGyARmg0VRn5rDoByD459V5DztQDOfKBxzQ/TmrYeQuUNXgkKupD6KZaX1AtGi1
TjDyxSukc95Mcxp2JjFRrSPeZw+E9NwmaPSudtdkk/k6bubeEZMMN13D2+2ZAXcn6t9DqSCc//r9
AXYSs2oJGYGHH/Ndp0zrKa7DX8rWbOHlWbmC7brQ56N9+G2XQYvmGM/PjV1hQa6PFZamIxgr4o1h
r8FkiRDUxOb5Sws+mH4nL9za+otagpGvrQZUNxB5BdpbqX1W8EjHUnHlIaz7NcInXqz8Pej+ud0F
tsrwWVq5DEOvisKqDkkZZThiajh6EcQeT5VEILjczurWkcR1m78B1Y1iV7CU5RuVX0XOhkpiitYD
DSyghSayyCUhdLd0flmu92d87qtIpJRSqoH2jZclXnnZDAYpvQUONe0QmiBQH2X96PutryXLJ0vP
iGnQ+w7sFs+KfkNkRzOI5Yt5PwahVDD6VP4sdqNIVCwyNnV/kCH+JHFUg2ww1lK6UOIZ9XsjDVAW
HYlUBEKC5cGOXPm8yUddFLM6WTYFgsYULO9hC5dYkDoynJ7CPr+j0Nvjz0OIJoJUydhMnYPKpFRC
jQFZPv+6cy75gLAnTKhX55KNLJR4LAp0Bggcxr0UGNrzwpb3yGxuAFABWy17W9tdCXCNzZ+jyD8n
spWhsD2+gzRlSs3FzM+z53nIMuTyrXrUUTIXfCKmL75NIDaojZRfOARYgwaaVotEfIoC3R/aG1qZ
QyMRbr/cqqYex/+aejwYkieEl6ocNRXPpe5FFHWsfTCcGQm9yNBqu9UkRP2R4iJownHvhzZh3eiy
jm9V+TotOJNoVe1zW9Lglc0Snw/AHRz7ehvT1Sy7yg4srerwdc34f7gKEaYYcKHmD6ORh/gSUlV0
ar/fLeE7UMu9Tpr/gjoO35BT/p+2In0uB9A5mtnOxuP19hsDBY1fHR6nNHiQQ4hZ5Ctqcwsjmrui
UdEg3CD/B94BFPGQQjTdLBsgHHHzaCLSWR1QeO5kt3ufRZRFU86JcG6662RWpCZlI/UDHD5lHoF8
GthlLlUcq0yAL6lp3murAO4XgnnymtPjcDD8+DiCZARLZRLSH278+7QajWGqndvyghCWS+hhzjDu
YvLWYyxQdt7B2E3DeI4sn6BsInQNvNFv1QBlQxeyWhtpU5H8C8eACqy6EzLMkb4SeKMEoEivmakf
IxKGA2AJKKQdqmF4fLdMSFYRW3auXOr7xTM0LX6VS9PWqui7/lX5Mx85RhC1g02yJZ1R8z9PYHhr
bP0OMGDC/cObbIFeOiFuL7HfGfrvNjHvzxJ4q0malRiSUIr5O+dzauHnIQlgg3ULwaGwkk/1cwA9
jL2hI9MMxBewPii69t3MjAAFmHxzHN9jK3GV18a/2XYlr8oPE7WHw+Vivnljo/kh/5NgjHROe+zW
uG7GsSXlIlEe8zGACGsvgzfMc8miQrcq9EAaKC+XJ6VY/dUQMycY4yJdrWFDeOigJSuMVnkEWjm9
jmSEdU9xvGdJgv7pvqIFGpWl1LrXBmsV4a3FhPYoo38RizMNE0ENHDgVeqAW36vTVlX8yxBSKGR6
AZOhLoAK98h20iDkwxrpxNlhFKYhqVkGg/8wonnW79HE5gZdJ2wf+CDagRlAt833/L/6voU+nw0P
Bgd/a2RftV+FiaPOO6WC2GzctkvSnGSYcRvlgchCeYgRNUthve87h54MIBCWkAGxhezfu36/IUIz
+dGJLU2iiDVwUxSheieMpGBnlt+LkIj2RMTPjAPmw2Qz5nzibevWhBpKUkxGx5HxN0cVi/mpQhbn
YgGnY5Zmp95S41pXyhHZv9NKIHspZMsLQqB/h/vlECoJQs83sBDyUqsIDWv/IxDQXhD3fvFF9OeL
u+k4Vwf1St6n9fMRK/s6TaVUzZnHtVZYcrLeuvHReBJl91t9lq0rEnK+/pTG4DcVrOOg86m2tW/V
1yNhGEC4dFuIJu4LbpvsyVEOXMvD45IJ6BQokQbaQ/1TuSGYnwbs4wZgogycgmcQsOu21SWzNsKS
6EfX4K4ZGq2tL3Jrsa7wu+0rcWoodiNyyjJdKxoZax32/vzNLGOxZWLHRuDDil8NTgFseZNpcKvt
dgJCUtG/djbLMLyV9i/8t3HJsyueKaM6HLjDiJvyOc43UZrds3VS2VR4jSvjwW/wHcLWuv3MYDh5
E1Qy+nmKkiC/jExNtnVE1yOrHUS19AKlkBatptb0yyeB5zwjQzuodWkO6BHVfuxHH1tTNrYyxUkc
0wN0c5m4zdZnpgA3vfGvIVJBk5djXisp9v/2QVwagmT973HEFjD9Wju6fjAiwiFwC8Kk3T5SKBeW
lcWkMXg7qmR6SeyEblY0dA+cKniZzV4wd6fQ2KreyTCWs0Nl9S8+2VJC2MnChx+rTrmWInWqsXLA
sSEYJI5dAGYuVQBi0+6H5hZIf6gGo/6HLdfJZqk2dJHR2laPYn4eY2xrvcstDDyC5gdpcTz4uoQ2
rF+RnfIQxreV8u1B3rTbenvco9nhP5WAfKRpjR3rq7ckUVwdopU4/I8MhWm7+GgijARkKRz6E5gj
rCk8NWx2AuCDAXf5/hWezaOTkId8UwHAn1eV24iHlrhc0IJiTsmlPC1xw/b1xvGpsap9VXHdO2+6
QGb9OVKiuVPjL39HDEw2aYDB4fGNbRwUTucmhChfRCQKxyeFt/cGHrw7xnXQgcDkfl/PDWN8yMSa
Usbsx4GSVq275oJ0B8zHaSa1JWj9hylz40OJckRnAgi3GvXMxkTAUNx5Oe3l2swCYhGh45AYScdh
Av7kK8IqkWB6bbklWFTXayFDCTWHQTp2RvRQ3MkAsZDej0RLM++M3X23MNOigjfY/qXnXRx+PNMn
MKLMBOlBh3yjfCbXx54eyH9FpMc7wrH4LOoW2Kua9Gi9a4KEqXZncMY8Y4MYpAkJQbI8K83EK1Bc
jv47R4YO8peVVpGUFk8YheOvAOQzUetCQxpZHY2G/gfcBEYtEMBpQ9NFR2pP/sqxxY3HcQ4wVMNe
ra2J2BYYjzf2A45O7jy8iYpY9Cpuuy7qWwBlMMzJNPb4N4waacyw2ApOLZhy1BsrBz3dbK0YgvRt
xNvMRFOPJXbnTpvXdJc9+S0Yj/CKm5AAd45y48VM93IPIsFZawiNGfIqGqjKXNc8mVa8SRcrdwIk
5rgzLmNqe/hIO/KQU6M2JxWzA462FRQK/aum0TBZxb/hAOXtODxZeqJ60bOW2Fbz30Qx4NA7iL7h
yi1EnwVhgmah7yTw9Xlz7CM23FK+P+P8Ml4r2ZrrDXQEzu8HhPra1jVdL3l2aC6oylf8rRo/yn5C
12fiwoHk2jhUwabuyDPHTamp4STU3DOX3OY3Y/7eY1Fvr9snq9vUZfjp6HkkqH55WH2k71zSnwe9
JqTfps/Dpds32EffQD2BznXf7CHr/zHiN5UCiPh0x5QgerMN/8IDZYE1ZJh+yG56W76j4FEWBM6N
ARFTSA/PuzfkivSFDc+9QYzbKTIQddQi4K/wukNi/5aTOhRyC/PdYTVzZbsgWp5MKmz02SiQzzwI
F6gsJ5Zm3aYdj33e0MZjVH24OQ+GW4JKqIBbWwajiWWdClUUdPBrZcIt8wqQERDYvCmWuf+T2Hv7
zMn0vGXdHfpMoqdRJuruXJxbvkMa+GFZsPB5Uuq1Ffh9uX1MqyRhvdJr7Y1E/M3bXIDeBWDzULqT
GW2XKSqhTZyg4NObh9p2IqELwWAcJHHUVkebXDZoarKJVbJwRWmM6RYCtOVUT5i0eQP4D7sB/HUb
xLaLXiQKYkx/RDwgpO/cp1LyG7VMfxT1FzG20lsBanvyjX5MZylny4Teu3UI8GEdUITkXmi87AUS
vhbTscdNsnxQub7iK7ELczj+Qu7kUF224joBny+RjxwKR7lUkXdZU986Pb83Gt9tvGkD3h3gjime
JUwK2v24BULnBNA0DRL/1dtQxUWZp55/5q400bHI0T4zI3I2r/lsfIc2i/MUd82/OBtZTj/9HF2N
OdYzerCDyaERzAJJQIRPzjhRdNSNpBIDEOUlYU1ljsu4EV09LIEObBRFzXHl9yu3gkaO0ZPjK/Px
cSRxIFe61IOEvKk9Dj0iXUZP31t1Quvfm9MSe80feP/gX8svwH9jAozMuvp0xsFjIc9X1ftd7xon
bN/L5y/0Uan42JehaX37k6RZFyy4S52wA07LZ8a9qochinMmXqPEM0CVHlwjp6kuhN1XFYkjN8MQ
zTdWTLfXx10Q2oqo3mHEOcY45gDjpIkEvbDLSm7yTY6BipwRq4ltbVUb1noZpp70rF54ZWlq0i8i
NO7ER2Pafntc5XCGsBZ8Y+ruapWkOdl0dlQ44x/Jzs7vaFYUV5tJ/ECjiYzjNC6E81q3RMVWrUwP
IBxtw8N9pvh59sSsDMGVmgCdmBtiBcFZnMUwg+5onmKKdX5OZtPgD04WFwWdWbs6AvUTJNjpE8fq
2mrFashL7vclrNEGf2F7S7Gaxy7Lvaa8pip4gcmQSUvRBzFfaUWNxA+zH8lmNDNyAU4HW4/WENKG
mT0YeBS17Xy91Smwuc1dank7ihsag30sF4Y4m4M8jvggou61ppEiSYY1v0Q5oWSFDJO/gy93rAuI
KVRTZkzio/FwxqnwuTwVHK/AxqU8E9vdzl7r5uQMRtXGiR9fr/1zJWjhCfTjrZixtsR76QILU4Jo
JMW/t+YOms6Mw2rS5rX2AAZ1VeMZIjXBbUWZTIdXpQCTvcVoRkmD70vleE20P14aHTy4iVRMzsZq
LhPk9tQgrHY7b6XBpcBcnDdOklWzvhp/wIVyDL73El4VevL8SDrZaCsXiLHr2FiwEIGq0ZrHpz5B
6iIW4ps/jxMuMrFMFMdeVNgBbDPekLxhxx0fY9A2nh/fM/10fT6dr1apCLucQMyId4qB8AVZR2DW
ECLfyLmD/tX3kCfXoPg8TMun+VhcTwTQwRPta4QSbVLMFocRIbixtLTt3FpmmevKPADQPOeTufmz
vIj6khHUkKXZBuooPWqoEioq8M424UfCfoFwdm9FDBFuU0HkuoV4DjGQF16tEotSgitagzstazL0
jAaCDD5oWXgwK7HBjJIZNsnUZ/C1IinQQjyhkAseaMFlJHP+Li7TodMM3SfXC8jMimVx8s7IEvZU
1eZZrEgZnklOn7q13VKg/qsQyThSC/Z9le6GM596z90uU8kY5QJiNvWnWlxzLkz2f9KzewvqM4Ji
S1oVod7eBw/gzI0baGA45nfU4JJOcP71fPbp+/rMe0nHckIkF7nLi/MWS4/V95IZt8qjOHTK+dqP
Vh2TUeXXkE9fe5LRQ3w+Nqbz+ufpvve0eu1NMt3MrS8rNnodAmtn5izbwmBYWXfTGqy4r7t+fAH9
OPuJ1AfVrYS1z0KDOEbcZk3Mnm/ljsuKf+5pfmEmKlrjpXFRsWOVfPxKii9R7bm6DMDEGHiOtcEw
O+lwoJfKvQ4NvSJPdc/MGJNZs5EmR6P2tuKQwGgirAXerySZGk1HO19+WUz5QPwEDFPnaJctLX6T
3e4SwH2nCgHNQa7+yD3/09JO/io9ImfXImfrgHHb6SqLjalSCLtxpgs4wDlVUe7yXhOax0lSAGfx
Rb8CJbCcWS+wg+Q4PLL5nMjdttPJl1JK6eHZeszTakTbzcedz7+HRaeV7XZLc9wOmCzcvv9vWSIx
Kdci8ppIP7l58IQ1r4qJ6QHFtfQAc63RbU4VoOXzWTatNu6nuQUNjp1ifiindEY2nNrI6xrqwbtc
YnZEROfGFtXBdc3lD5R8GweU03Orl4SIut2H13ow1vBfMqkX3mBSw5pp9S08GafQddB40cQbMpCR
ai6qTz0FFjalTwIlKE4G43lPR9Nxu1m9cze+KelcAJ5TetXsgD+yIfxrPsn752VcKoDFV4CkDuXk
TjfAh/iapBgPMAiKjMnnpFVuEA0aAykpBtCW+LWBTXiqBer+RSOeKUiR87Wc87u74G00B1f7jfjE
0gdYmQyCJkp92rC8giG+1c2pB7TJm0TVWHLSwIX8lTFXSJLiRFsG5ZXh3MAaVab9fN9maj10xmFP
ePmYUWVJmwn4nXV2dYy+H+oJ9upL4dR4tukfvJmOSlOQnPIu1xjs8jMDhLsNsnR0oJP+iiB3H28M
5QeRxDboEJughxMqa9iuTHFAhXU8S0P2T8O+BD0vd07OaZ+5JO1QqJK4q8w8pBFDA2m1e3YBJNEJ
L5plHs5U6zeVe7x20dnC+8BMcJwjwEdxBbFV7FPK6GjXJ+Qldc/S9dQ/wceWQMdGWVFTdMkCzJ9g
/D2xdsgCWeLmMNeAxCByXkFyp5ZtmTkJ9VIbfVCqu/8IUhMWwKCAEnuG3gl0TYNLMSvNACbTuzOQ
23n+d2Z+EAU2Ox+7zaxhsm5BmG2MhOYr+I231lyG99wixXs6r3jSDwaecpKhLkmtBlEowZyhke+h
FgLnFjKElFX2LxsAVMhA86Ge4JWdndqBDOG0a7DGXR4lL5fAhoaSseQPsNsVq/JPJMoIYb9rlE70
UBHpffX9M/v7/T1hEeevp4q2hPh1aN8mAP3erIi3PhRjbxMsB89xpfSGaIOwv3ClXAt1h87WufXe
64P618DSp+cHw7DE4C+rnYxSBJde03cDHAtuOlcHBxOhppwVhG+Wlzmq6z8/XCaMwYlb8xi62HBf
4L/CfuiXc3GuemLVy9Sn2AS7avYTCJseBFeAPT9KEx8vEF9Plp2kVYtpmcMe/VkD7byePTGnNoSF
woprkqUvVzov9UoQRFU5/kKcqCDSvVF7m5HR3ioCd3xVjpGd2NteWLoJM90zx6eYqhb3cmYvv3m+
Yp1seliCgpgJGlDpcTAHWu1ETWn8xnGHPN88tElPN4PxT2qlw6hXYz/Wwv8OsY+2cTIxu8PhQj35
T9hgLEXVI6zAV5qXMYiB1vIDUrrR3BTRWtZmJ66hjRqmbB18Wx6mZa4I7a3fx5vgSiNeNCezw9Fl
iMX2YeNgSICf/MCd/Dm5Fuk2zMuEs2T9lMnzIUdF2GdACwdvyLZuhRpO5mWcd8krk4mXEXmlc8ef
2hmpmb4sPPXIgk6VccF/DJr5RC6MpuTAkysZRNipWgg8VmNZVyAsaGisAnFxKKEXPpYvt8c/2Mb4
D8AMeEvk09ds4FqBGNq86jTWZLaoKyHhpU2mj0JZsMTVaePG8La5eYhE3ZfG3Q358duratalMeUx
NxM0f1cn2bgx21ADivV0jEgQBKKPMaZe9BdO/5V0/F7+RxQpwoPobKKX1fj3dIN7u5u2pYzuVa1C
KPWge3VkrA9IrBa3bC+zJVCpLtEBW1KxMfs2JGzgzEOoMPKtKrK+Fa0zJaOFgoMDqf+8KcLmdS2v
v0X52losbLrnXLrzQxpoRcGZqrdZ28QsOVFXdRXSVCbUMZZ68hH/cy0zcaYTAHaoqSMyuqlMIayo
kbsvIhnt6UDLYPX4EXtQbMTL0v0qKvZiT/UXPwsdrqi8KYvoXX3gPj2mt5CCiEPEopPRFLGAyCc3
ohV/CbcfYuVHmetR9+qjAlUVccMCBEE6F1hWlnQjNWWjVpcMN+7lGJOZ5rpyyUE01aLfPJYuFjKM
OF3g4og9aR+w+yLTfocFCmuTLQHUqJIq8V/OWx6Vw9LCBZ1woo+0jvsvzbVe5lHK+Dps/U5bFf09
0oO1WoVYUMiVa6znuNHZj42zWVf/4meGCGnh+Z3Rdl9mhD4g3IUfanRId+o8C601og7P63vrJxOu
R79ABbuDnqivODyuSC0mCDjV7KeEia3KLx2Q+RJI8pm61hhFSB2oq7CTQGSEDsZ9P9eHK1ZgVgaO
aMWRC+eIdK3xqlMU4UTAp65IiA8XG/gyEFlVRtu4aM7kIQPJX8aTDo17KEQOxtC1SYj8Z2Lt/kbG
CBs9t2FhqQvni4816yZ1EQaLP279kKJOkDN6iPuYWCGNdCuesVXyW9qOH116CfSucc801UUE3SNa
0ibLyx4ijbFkBdwy0MXmOjs0nOHhn8f6H1Cakv8+jjscovXJYLEsa0cbeMvzYpcQVNtRdVeMVJRF
HNmlBZLdKbej3LJRWk/mj76NDJO+sMkqVrcHhfOmB7a/B0S+WcK4Z5kgdniY1OgQrCjtKgS1x5Re
5EQOndeguCKuguBYN6ji1Vpz4SiUp5vtPm+1hw0Jw0CS56KpYMlbH0oI1fmyRnidTH7hObkne7MI
PGN6I7P83RpEdCKJdnBwh/Cc7TG3bD9XfPxPVj9l/6JiWXB8PMPYeT9GHz0U723VfprGoIfxNLh4
TWCFS3C3fauspU+viy5MLnYm0gfuVqKxuSSB5GOxELMrbHM8/VZxN0kOK8p5s4wFmcHEksuNkUcf
krTVdHfASnqj910ziIwOeQrdpHRuXA9lWCeG0GpbfJoKpLlkQKR/p8vW7NeqzWMyKpqx1APIG27R
NKxTRmS+zn+jDwKGy1tLHYbioCYzN4xKnYi7TvZHeZbmxBfIveU+qN1MxhUZa8mZoBhq8QkJPX8f
EAV+FdfeTrZxrhS2mLMpLBxDsm2Yu3CsV7DCr3PIR/2GIajuhQuKKeR3zO9dRa//tbkWzuZvFkmR
/d6mqFkKBClPvgFuSIdFA5pCr3A6MJMoAI062xS0aHN0j/erRjo68ByygwllQRJMRkFFLNKqoWW3
Vzy0bEm23b3IBYHCws1n0oXiwQIEsEQ55ji5EYz1kuzR/w+xlVQQqQtg0ZmAQq3Izc1UiNMPV00m
SWtSFk5fJ5k8n9RHJszbLFoHtmasC1B98R53IsS9592WEV4pJdXR6f3rIOgWkijm9OVoMuoE2xZ0
bsfneyr79SVaYm3bbIjhejFpOweKhWP/ODRN60Zu3+BWXbJxRbb5sCNp5NGCa1Du6TYfaixULTyZ
5bIF1QeXX7BhK4XXcUWbrsjSxQgQfSfiuhWRhXQRTDQRCOqi4wpE0LLg/r8ZFESU4ISAuvaz4usu
tTWsrR6qmEb5UUKJAOwtrFYp89B/1LZxO5kcrdjeICAXBEWBH1/uIVzQWOY5JEx8AJ77NRkifneS
FOqkO/4XonuS0SR7TSnaVSiqCkrMJRw2MrQrlR+1W2N4h8fLOpI3PMDnim3ec5bp9z1G5e0M8W27
+JD0WYxEr0R+3+ejLKn3Kvj8Xz2e6EcbXgB9LIGua7OC1CBql8ONPzARLYVkw0MM+0dKethuTyuP
6y4WxUtzkqntoQTLX38RMjU2jgi5o+beUfaUNXZE2X8ct01IC64S17CRk4qV936KVEqifJbB2kdV
frRkp3gWGKSCv6cJdnRDI41t3OgrFsrUN/RmIEBzMHakUde1Q2kI6472aT3YCrLh3vyXeA7H1hOd
QiiZ/A4GmAYqPQtxlcnsBO/uS+D3qW3rRtW8yNDhLERW5Ay9dBihu8/taPiQOc6g8QLmAaiNOSAo
VDHDkAdUriHW4/bhDVx5IFQGj/rf6EPnVlIeV7BTfUhnX6C3Z2mTxlRqeSKiXdLjxTsG+4fZTRI1
xIFKAbW1J6N5KOh5gZghTfjS5S6Zt16WvpWDj9NkgrKZWRC2xNYcFG4BJBmwF6duhS/z1RX2XNfF
vVas+ahFc0TVHW89ks6JGMeZzWCyh+9EsLXbd38G3lMGI5qnZdtxaRR2U6r/dkzcsSY64xMFxxgx
vGsxa6hDZXXHrxtJnx5na3LmGn+iuH8p7uHtYzruKjnE56aG6NvgdsOW1eMTgGt1WLafeaoxJxpi
4vpHs3qM/Dd+JKkVJH0HAJne/IVxrR1QKYGcI2IW+olsBH9Kc9IZqrW3gB0+FYov0fsjQ9cgwVLA
5OCiLvYPIWCOkcRWOB6oWGFTJq7URmjAZ6bChjnpoktyPlaoZsSuAx0AmO2erY/kpOwvoHibxAl1
UD4bXx30LpMUhb+r0wslQ7utZ/Sx9lhflrtKg1a3ZjN5EU1n2+Zs7QqWTa3Ln1RtT/OQCZFTeO/d
mIDiw9pBVb2lD94srp0bMmnQPoiuiW6hflXE2tkUhdaSk8VaqSVOywJp/ISBX9D1xPVVeYdMaxJ6
DI3vHH3dglyxNAs3uRbylM1gr6sKcH5pQmTIUJhRsDVidNotJLrLxx6yoLDanB18A34PhfNVAHKI
1M4M3rRRnuxgB6vl48UzTu0vcDz6oa5GDJLoZf6qaLAR0IegE+vixFCzGLJelrdRTTZoS4rI25WY
2RZIPCeClQzKrtzvvA/1PM93VEAr1FVdq+KrtaTjU2qzfc8rv/Yl5HHVPmZIsEC46VbaCoDIjENF
O4p463bqaVLBUYb47c95WV6u3+BuLngNBaG2mgVWQhV1qESaaFliYPavJ9DsnLKxUfaXvr6RaUBF
7ij3UGMPQ8Q/EPbhJvvlH7OYv5xEm2QrvMziNGOADSZ9a5h41e6CLUnajMHLRA66K8Vu819cuUPR
5jBgI8tPdADkgV1wNVK+7QfADH1x+lOBv/HIhiK5simhKH/AYupVUhWgq8dnJnEMm2pSDcEAed36
DJ4jCS+ZI8fa0B/MkmBVbxJOTwpUYJ0UgfH7OQuPa4Rns3Dn/14BdX3Cg2wXlo23KvesPV2K1TwZ
Mirnd6riL1SKKEFTDmVYFBirNPTkDwfFfre7w9hJpUTuT8tqvmbiL5awBOjlpVaQGT9Q/FQ+utKF
N+XwyglntxcmDd/GjXUYHcfjdCqetI4wUECeDOmbBwyLvuEqcaqOMK3AtdkEwju9BGjEuFX3Vpaw
9NFXO1k0Mw6JPNpCf+ktO84CvSImrlMNv2to8QVUrFiSRxmK8qctZo3qqWkLgJ42b+TLB/NlS/CW
Fia1kfuzV/F115GDGVEgNO7zh+hQD7nVARtOsQ42V/WG7GNXPMkoTqxqljxlkZKwJRDCj+aHOlTS
WBeG/s4vk4838pZ78bQXqkzhZ541SkqrSwDLzaXsmIH7U3uper9tiVFYyN7gj6Wui7U7yZmQvXVy
CChTlN8cvaQJBR1JbnVJBR3l46FuEHumKfv5epYnunrOvqH1pBY1eEs2PAZuAswe6SjkD8+PP47e
mtLjh5bDFG9d5+jvlNjY6qOf+QPtoAxUBVSR0iaf+6+7mNGsJ3PUDvA/jeSzu2PIValeHZO4mVX3
Xx4bl5R+TC3qzx4EHvduaMa6ga6eAJuKxwiv9JRGKhs8XD1h6nfgWvFzSSAFPPT9W6xAPbFDGyTC
zxdFEV6KAClwftKXII20HYpt9J42l06JfSfErzRCIQXjMchfuZXl/5K/ZsopYXADD39frIiPCNpr
p+vIIeRnBQeYkDz+HkhmPq2MxlZqm9Gs200xu3Xrl8F5e2kHijIJPyGpccSrjjVunfvr6Ugaq1g0
bTW1fRE0IRXXDOssqSlSx+PVRdfN2yMRMkBVUro8lIqonPMdgGqJZkf6BxwRmynCedbBNlUGGLvv
6cTkR/CVdI3LQUda6zTwGsYhk9fo0/czoe29A7fgxZWRxgRZgC5UeLl27dMisoewkfyVxV5dDuDE
k5/ZVkZDRIt+M4m07x9CoDaxF2927EFyvRs4Kk1raphUoG9HYQqOwuEbsKoae8UDvpRWhqshHezD
2jPJCXMfe9kj4wZlw4+dwxgOeTBmMtTyYCFm1sa5AB+XP2oZHBsopX5rxmOXBWsV5a1x7vueIykQ
ZQQvbXB1Pn3anR74plbSb8xW9hKtjP4FQFAmVDerS3IzuXPheZ+huww5oLOrCKTznFYBe6mCcuED
LV6jeKAC2f55bu4iJ2i97LU1OtvONcaBKzOeiAZQyvJzOn4OvZ/oYyx42YOl1HvrdAEFS1r3y66x
uyJm1z9Y8iMc0UGOENAmcNIuciJPhVX8kF3EkgTm7prk4YWT6f/WDEhcHiX8xLEqGjKyocsnpQkF
/RneiyTijruBKVZyb6udNk1UO18yAQKgbxrZaCcZfokRKLqQszJweYGDciVFeXAXWeQPkubrEqSj
ScmkGizFQMOgMtL3oUldeD5yHveAnHinWbtxTuo5U9paexj2peLaHb/Npj15NsswuNRWeoRfpQLL
QfjzJREidnz8pgmlrHhk6Rq69l1soKJZwC4i4oADzCPYb4zH93nwV108ZXJ5bLqzjJlDf6Rwu2g5
VH9MazLYqL9jw6JSBo5rQXe4E5Ajdqgw8TpO0W+hHRUG5SHDHk7aC8Q07cGf+dFYyowEkZQti7CZ
fm99Kc5TbCxWDB9oreuzPo3480ogR55SF49nGMmV6N7UuaFy+9bfcL6unqhqsQbXVZF6MKLoRNcj
g0FWWhLLLyXNhqVT4pi7o/m9eW287AcaPuwncuoauVmeKmrcsjHjl1NiAXolKZVIQnPvmn7wMWSL
0W4f2LFIkz+BGYtdOQEVUk56ZPkrN65g1j9bLQbXEamtziQBB5VmR0fK02zpIZk9CQlPMEd7sYaN
qJja2VqalXzt8buQwj+1EcxsPSGwQaLivaovd4hj5jsoaCvXRu2XlHAw6cYkBtUGcCOIuXedzvtt
lMajKGwMUY+wtHgn1eEmi6ZfZ6Sv5qpMWfoET6kwEdZAn/p20swrq6uOQEky+BW7Q61nvJIP9r/s
YeUY0px3iU6ZB/3qXPczT0VYASexmeny+X7CwlcZ2td6dPU2t+A7UQe1rsa3n1JNHD2Wk5I8trsi
4wmWCRpQh7VwHeo1WvyzI39JtxVBEtWAXERb6I88NsC5ybf11xBJnM3jBRzdJZcyj6DqJf4tWQA1
KC4oEou7DkfOPC2KdtdEK/i8bzOTOtLnyrNA18JsC0gGQ4wTN5yd8nZuy4niQR7+KxKd1gzc4bPr
3z63GekOwJ080VpQcUXUi0GGjmbc2gdclpCMnNs0TZNSSyOkyvONkuZWUpHPhjYR0tRTKv0dbh9z
cl5Vx243OsfMaGsZPrP+2KEXZDYz7rTwlHCt1/Z/w1vwGeFiKPCd+Jgab3S4Tn7/XBnpqX10i9Pd
5zu6Aqw8LAIXy4umbiiJ0uPwnwj3Ok0FLiw4Uw3hyUlBB2Q+7msSPMAIxLNy5pBbjhdGnqOI53Hn
meroFEbYIevMjD5V3RUaOxsXI5QOvHGgGuD7D+19TlH3o4cJMmt61Ic+Feu9x1+yeRFwA0IFuB9P
0gCmSy9hF4A1Ah+uueL+G+jDQezJzpFoh8T+G+UjmeWhBiRyQTuAm3s1htUFC/1tTEYpkYYWzLVg
Y+qJgNJFuNqjYsINrF8p1lbgJEqCETd4B+AuZaahIetAngcSgPYdtca9hk+0xzLYBC45fe7o0V5l
yJ0uX43R3Z1LZjmsuqejuUw9zga6Uo4Kd2Od0IFGB4Tsw+5e45v+PPfM50rfEsHvw+ThG8QSrdfl
4KYKKCWBXMrq3qD2G5DeEkKXbaxVSBzLmra/RnweF58v8ZDGzfdL4qRX3ekVQGqTiAQ5PN80508u
Xd82w8M/p0T4DcOX/ouJQShsMFX1Y7NgQlaTtexU3Tg3+u4EvjuP380sypATxS1toEyZXeYPPKHi
cW+Rj417WgiO0+PngFNb+MoGuWwAfXIRMA1sNUQjol2OcTGPsz6WwsYGY7T5CXBsIoEu78JwzRDS
sw8xjCGHd51SSYh+RfLX0WVL4CJm5TsICxC5mfcf+XY9lYGybVIxTSWCwyJLuMUz4ImkqHRyj77k
uIlmyyfz2qB0p13DnRaAynBjdNpukSEkR9UZ6R+b4Z80i/awCSCmhuzCofkHiGbRwTlaM/JilcCF
jGdD4qCbU9Un8kd31yzAajCGUJBhfSnGtMUunzQ9iU8Xwtue2zYVqnRnN6gQBGFCNwL7ip6juUnW
SgAvFifA2oLrScghXqkw4IEon3pTSXI74S6mediyXiYQ0YRxriVUFW2POcHYvLf0j8mGNd/Z9Phq
/8BkA8XuzjQQnM0iDzvC1JuMiJ8e6pHU7bv/HA8EsXCG9H/8cn4luyPNoE1zJSE9d3qaMBjmGkdd
36t6tk0MOEiapi94jHB3UpHa0k+LdaqrAn9PPVEaA1QM6+sA5bOQRBkM5Tk/mDIyB3XB12J5PqNF
ECZx6mB95cDcfAyVF2rG7FsrwRXbsu3yVXHVKkf8BBqYpfDdt+JjPFGq6CtIt1dEHWrLK6lRColp
k1s1kqJ4PciX3dtYrCOGGXv3cHBIjHdOffsy8oQiZYW73HrlXaH5CAo+PLz5aEUvlcXcO3qWN2CO
ATHl3KGxp0Pbuea6axlsYOtzoTtsFlZKdhaMDFJ1EMS8ItuY/tJqvw4GAVZ1JDfR/Vd5XEzd2P2f
Tcdu51bURDOWYDDzipgerPhUHJjUj4vXYtBp/ZDOiytSITytlR++fUX2wk1FT8rV9CGpzOs50Tx4
8M6+1pifeP/vYVSr8kTIXepYo8dzjF0sVQZ53MJgGBK/MfY20jKtsYolTaI/dS2fhqoza9QONHbU
6Qvp3PFFwAJsilS+yT5UjeJlMJJXIMshochzVelTmO9vPxbMWnACW9ih7hPkaZpKEhvT/TH4A+vA
N5KPbrnxFe4IHdj3GwDveQ+6GB8du79eTaXAt7SrcJ1JewFIUbsNZePCOEubIQb/58yh5FNknQdW
/I85hHCcQCcRrfM4aG3IelcHnO6Z/wmy5OMhKj7/1slhZsXwTuzKO2RaX3mw4Ohz6TQYVQBp/nWS
clcAFxqZAxjoajMCUbmAHwC9VokVU725koTCRwu02h5xLyZ7c/vD65XqkVGd0E8CLvDidRodC+mk
CkHpIuSnV9n1/fYTiqBWQZq7ewuXQZQqqqj02tSdstBW/nqaSL/wew/jrMIyrz1jrVvtrxdK4D85
u2YJm6gHcH++LQJk/vxh4Uy2KwCaLaXOsZMc3pFNa+W3oXXo4G9TczfaGqWCUJVUTFaidSJXIsWJ
p9lVZ0Ia5Acs2ltPtRHkmOoYuyBm7NHLBkKI3/fiWOC/Ih25YD5b9coQ74MeQEc8Np/+0p547k1m
PPKM7qOPmsQjI9eNnbhqByG2fy+bFNTh6mpoN9jkr9tlKWchfLmKOrEBDlgNNDF4zM5KuOnZ4ZJb
EaEKvEGG9RpiEOFb1HVF6norj2AyukI+IrnT4ahI/Ya4GwrGPz+yLzJ56aVb75ydJ7sn+jPG1D85
9G39041rDQGK+mzwkfKr0hGsvLkWXqxIr0idYcZxBheKOd1l7AfrrNjORk3bEBXRhGGRN7p6IT/t
Ac70MlW4qoWyNEsBxJiqpIXVeUK/LcvLd9pC2kST2/QyRTzJ07B0ZcxHKeaubByUiVaFcT9aghXk
fHm8pz9Dwctir5uVG/OoZ0mhN233Et3bDpRQ2jP+gusUbJ1CrEK6laVjiUNcQVrile03Tg1U45ip
MJcPGNeo54YaXJqMly17TuADPM2eGXUuD+h+kuHSIXZK+yKGFFj2d5RWc6IECoWz8RmwtAso5/pz
d4GIKc4pJacAH0fiYS47/qDQvYWfTnX3Yspb1ivyeKd/25XHX8yVRAnguRVQZdR1z26LP0V0XZsA
9zb2WLkzIB0vldK1QAGqpGXYLy0okzR0WGEr0nqveTg8vZ9jkGsuQ6wCdwDB6O0PifXcyX6cacqr
WycLBoY8mn8PQN6oJEFONZE16nCg8SIWmfQ2ERCUvlvaDMiBtH5Uj1h+NMaBHg2hb8EMq1RMOZbs
ValxvolZKN0MIHZq47bfFXJzHj15TKMZcMI7kG5B1XZawZa4i9QQ94ZEVwPbkEfiumDx0CCEWjn/
NSO5ppuJvRAMnPA5R0QbwKaU1ONvzvKlLIKQLSJSAEZ6Q0KHe92YaiufKNTTK9lZvTYUfcPXxt6v
oYJOdVQcKW/bQFQTGw9uc65hG1INo917TfFrijf0HlSZMgUkeg0qjG2Czb7cCJCCLQJdX/H71QSp
zntV4Luf78jKwUNMm7upBbLx2EUZEdR6zCcMZAqh5ksbH2avYryg5vwc7+IvBRg8FSgav0UKStNj
J/x2QUXFpdXl9KeVNUSYVPeVftdor5TNtqmAnXUAM05QDxRAuyinEApTVimTlM5PkWKZFC11xi2z
RRYQ1ARnyxBI/FV3wcZ5yZen1WIFE2ezHbfBD+IgyNmJuLXFqGgmL69VSvuT0x6gVsXZnf6Ckr/b
JlbpD5RxMhrR6CBtmbNo+iUmasBYRdd6z2vMMuN5M4yxhGZTp8zU7ZdG8cmnENLr6C0M9DWq/KlF
eTPIp25OeApAuhwBWlolLFIcFWrz19TiLr1MsxjVsbDGT4ce7TWEhKrplRLa+yZI6TM0cV9Uckdb
5lzlARa05ElExsE2QqcgM3laTrlioY33mfqteVWxgO4jAjwSE8DxkL6pOs26KjZwXqOOtstdSqyN
4371HFrk16bSiZdmpQBYKJvr7tWd544Dz5QcVdbUJp9nEXix7ZJHfb87fWRV3JjqdU/NjESzjUGS
ijnuPKRAwPyz3GBPg3B1AK1HdIlF6cLZZzi+YNvl5ohfv3mVZ03O0q+sgWWfiwi2tpdH9naKOmAS
G/LmbB/P7Fy62pRI3jvYHI8bDJjntYqvgO0fO0bYR7/+3MWIbj2mvDUgKpiBdxp4CVg/hXPHMH7h
mxrHawn+Xm6TGQJGxYWy5J7iNpJMWyrlCGjBoPBHptyftlRgal8LSDxVtCG6bwt0xItufMu+MSGT
XfiPwGv8R9lRORABE9KxSmsFB45G+D8urQWJIuCHzsteFuR5LYZFTiZzS1t2tSLObnL/ddbDmtq9
FvXu1N64Md9ojHUB1wg+BcplkBUlH/oH+CL2R7tU68rbR4b8Yu8N3Iyr9LgRLxA0qBElRfxqDFhm
LSU+SrGmaxHd4Fc99lTLEcLceWhYPD4TvQie/jmDdWOHxyDNtjKZiW0UiWs4UmIfVw5t5Yjet+on
xTBHM1th4H9S6JZnuvF8mW66G9q16GP3qOeOipnflPASYKxNywJ1FbzK8+PVJOW++ydR1kz4rQZU
CS26kzJH7OIIR2PKU2SO56u4p1qdJU3owYyOKHNR6Qh+0lA8WlxgfwGTEqQLUXRfxModAuci005f
J/x8/7uy8wk4na+K9K0K+UKQSE2RJe5HKumNAVHIS0SjRzeBmsfAFcCxivTFHZgpIEoXoD+B53wU
pR41ljrUjVLYJOY7pdfh6jSaHKsvdRSbGjz9duRfvucetjinxjg1y1rZLBYdaAKgUGFc2tKe0POw
bxvRGZnNVfyZ7N7M0RMtXbE9cj/iICBibU7kC5ZhW53+hw+oXkwJqJWTGUVY+OA66bUiFHI2vvxy
gTEcQoW/2oYOsyX8otXi8wg8IzgQv/6e/Bagve6eK/9G8BimGNtoe6R6ciBu3p23TdC5BA4etQXR
d01Jrwaffef0NMxcOvNJXj93jCd+V4l69s3WW8XuOgTZ5HldlGT8TORDAW5ckgnDW2VpzWYIFQJ2
QI7C6ihGplWc0K+u2YPyuGZtlHf68lgVr7ztzodr96jG2CWWs78ERE5t1gqwwx7C/YwMlx1dQdKu
El12xljbGMB8/TtNiIfSjsxZdxeayZnViUfKqhGVMAfeH0ep8c5qXj6Vc4bmQ550l4muhgviapkn
nDKWbq8ObLMbY0mo0IYBweDT95jstYfZNi+RarGA7IQVNoST1xw57ooRsINVL3fGnJ+AhZis0YpH
7Jq9jJhJ1+OzRl0CHYTScolQbqCcGrsNgmO841jwNt3xt4uGW7+8L7iInP8iV1f6OIp3b8eoS0lv
taz7iM9raWfMhO205Muysshl0LjpzCer/whL6VO40kr/Kxzexu2iNjxiLzq0xbZWvCZXz+mde1Iy
7NrGIIaK9a5fsjDmj37oB1Mr4L6S9GM7jhw5fSAJGgcDjivOXfQnxgGfqjjzrRe3HJnmB295bFOZ
ALwcHXLjH9NWWEE0yuFTe8JCBntaNlMeOMARDCQhGBxus23BSl0mhW6X9awrvgzDKvl7Z4dZ9zv2
Qko0nsWz6H3okLJO4DsKzUyTQWKCP4diQlA53GIigB0KlMTEZvvokSZCbkUIV7Wq7+0fw2o+1MKJ
EpUtGWJZE8eu0PVtoXHfB9u2+9exM9g1NY0bh1vznKbD3ZZXTiYegTw3GUWgi9BNgLBthqgW04s3
6SkW05qMBAn/JmzDm+r+FX4U434WVNBsqhbBzJPOlNx8Vw42xuvIC6lmXXwvpztt07SBqNe+FsDN
q/4sfUBxl8vferXelmhi6IeV1sEbE2b4HTtWiT/UFJf5tUdur9jCTfcoFTSGcLy8TDWI2zFBJZJC
BUM41zK5cv53rUaymSFSVIYugsDoo99Y0zKan8zz3wu9oL+1DUPiCT+/D8emut/fU8y+xcXBx/jr
SENm/wL4dlxdFT83P2wkLnSwNuwOr07LW3LfXX8Wd1PNOpWpZQ9tyN3ywN/Kro7+Mz0pulLm/j9H
gcpsm/Uohp3lbqcmUDYgXwewSypWJYdntGj+rwwjspRxOAr0lamYj542kAdnoZ8cW+f2g1HhxXo5
JLUJbzz1tEdXURXHaUIJWCNHuHL+0OQtsWcJfbSjASD1+Csm0n8+v3xX1yNyFxgN1QLPAIIC89bH
dvkQYqsMpTMfZbdTnO8iyb+2g/kS3UmOfq9F3US6H/2fIyG4LlLjEltN+ki5N5Uss0KhbSUo0/eB
VFFm+YDOLDm0T2PYQBM734BDgk/ETNPiibJJLcUyRTBcfRn1qcCaQ3rtqKWr9gOvHhJPfD0bFtCM
rTbFs2GVoiXSnquOu7g/Tk5hOWwpjyD7NTlOMVCe1WKoynYeaPX5hc/ikkKYmpAu3hbyKaTMDsYM
6HQu6waCImRdwrkVTjl3uZXHcsDwAwbLFfuvTCYa1OwkRvvLCMMtTZW+QvNcMpT+E7Iun568iNMu
pGuImgCDrN3pokQUY/We4vpnah9oTM61z/E4sojDJ1kIwCrFk3Y4pBcp0sxV9BXzZweAIpq4PJjW
Uq7Nn3sc4lwZfeAvUOMGaAVTUvHrEMDYQXj/e8PLh7ctiBhcuSA/PkJ47vKXCAzbgqKm9XBNkuTd
RnZs9cJNHZYB7chy9BXii22azBhA6XOYrjuMJRox1wXk+p5ws03L3TUQyKvn+1HV1sqtteqmNvc9
4W6i2QyPcku1d8OwMCicdHrqK4lZLQ2SXaA4olkXj0w8V2BY+tSfm/XY2Np8lSumVSmsr4QwsRLT
qi0o3Fv9Jnt2pQJ0xIreYLclDHeAq+YjpiQbnWo3KUNTlMLXHoaF7xxhWeq/H+kZAq2F8GS0V0Cz
kHcvKZ9MdMm/ESUJV9ncjZMbLdQloR8TQ+mUMvP/SQHrM5ijMM6PIDTWJbZqdIt9vL1Z6QzHVRxV
ocgnzCPqaSRpNp35aDXt7LiXTjrfm2qV8xbBNHA4yX2a/1/r/p1gNPPepm8h49zP3mSbYqCJFVEi
QeyC60QuCpwaOX5svTziaUVv/lDDTQifigg3V0pwfeQYfO2mOLSHhVj4nRJi6OkHrc4qLkWes0aN
rE7VTvukTrMT/rR4xFWk1pAul8yhAErD1gzo+bGVFnHaiHYrAYIbVnhHjdDjLKL84hVsU7GCPWWL
Yx+1vhPmqePQaliK1Sx6I/cTPHH4iVO6sELkYxe1Dp6i3rMAZFTcU7C3fIiPZk+wkX49E03nhB++
v0C3Ki/Djqz64bFmniNQYHD4vvQnatbqLRihZzXmv7R3fr0XBcp1mnhqoBJlH87Qligwtd6M0HvD
byNUZ1STlUAkHeMHKW4IWUrBjeYhvWlSRTDXKs2c7WgGfyRqo+xCPcKH+r7DDjA63GcbsGDMM8zm
0m5lDTdHh9VEzbqghQM8NoIRWbA5hCB/79Tzq63JOG/GhvY9oss04a5rAHUzScBWSW8ozrIENVfV
ezI26pak7ozs5XQfP/70GrR80oN5nU1YOZB+ePVOqnT7vI5PNm8f7GjSni97zDsiZy0IjBdmRhtS
6vxGmkznTTXT17hbkfuYhBvUH8SnSMFzFl9dguGSlgsYktUZnc8ytxDV64OAlndReTjd2tZkn+t+
AExwWehMhSn+QwqGLm00MKEpr0xcXpNOsvmvUy7Q+E0vdOz4cUu9i4RHeUiB/4fj+xYT6Zs2we4w
dB7YIE7KoLc7ok+u3d90C5k9Xwzc2EJ7zW/IAGK1316CguqbyczGTtL6Q0GxIfcFFoU2mEz8phxI
IG+uJKcm4joypzvM5Z9xTeXSxN0lu6sc/UUC3Wr98W+ya9aT+PHXzIveicdcvqw747wNjaTmPlMe
5DQCyfSD1FEJ+8myNbkLK45Ya8EgqxP4gd6aMNqyYFEJAoLhNRl82v1WnI9WTF4aL52MXdBTLflc
HalbtsSZGX2ysrsr30pMeaKkWGum3DvjofHpv7c+xPYMW8XZZpw3v3JnbeSKK/aYggUlNLLgoUT8
bAkHxXbnTQqOoqZ+fdNO1TtccuVIuKAoliptaQqWekN2LUVdaKoZK8QIzYdAZJ9kXYLu7WzOUxwV
AXbtOH5tX62q5JWEHJkYQdRBWOpJFcEMJ6pqwg9d8sD7O9zn+BTGqeOxzRi5mGsNY5hMuBZE0utN
Ne7OkMLzxt/OH+gMvVfTv64PI0WXGvgaDp0fs0wdwnUnC3EbBuyP3zzthdMiyNC1BKenG0BwOHXB
nBaT5BdT09scFr/EDte38t9tmq0uscaXMjaakXBs6lnmUDm3WJrR8cVOIFMIqZQvG+99eYgu58Kg
uZB6FlhWEIsI0LJMRoRDEsdixlcqQI8RM3AT0cSAxi8DALnF8epYMHRHqGov9UMTJN4lAT4Aa5cv
dfcGzL9Nu3EaKLTQwz6s1j1aAb/8U2TaEsKP+Alz/Gx3kmX8HrhPDxCjyGOlCugQZgWED8pWaFPn
syeglR/WDzjuUNy7INQAkegGKp2UqjJ++79HxX17q5BgqkPvOeEGnAfwUQ0ZCoBCp/ljcabsFVTF
fbBOa/FoFlIKsftG/gzHFAxoNUQ4x5J1iNCNADaS7XEvdABVoqMbglRAtF+37TNWM8rEcKcb4uVW
cijWH9pctlqQwaTXvKEoVIoljADvnmYak4wsbL0gZRcUgkMO/e8N2rxuBxtOTg7/iJHFO5PaS5pL
FD/r/SdACgifWyX964idOxtfFHfifwQ9nHlMMSn9ECqMsIt+uyQ3hVLqkWYDGtZzODGUm9eMry0U
k1kp/zEHDyHRJZeJ6v2l/egNZGBWq9ue3OMTS7Q7+2jGkifDgS2tFlDHQD1Xc068dfUxwUSIQ/78
LQpDMhi5dAh6T4xXipLqWSmjcVnsqFZHxgYeJAzU9jBcc9mkrmRdauPX88ivHtezehpkpBwbS7oV
bbFEQ0BJUn7HhzyyH54ipy0EzK61KIl/f6i/2tmKmm1Xmfxi0ukvKOKs7USp3d8xJtY667pSux7Z
XJNWe3YISgpNqrLL//IkXMWHZudyCGooLrWyV1ZYBL5sP4wtE4Z6lxTvoQjt1s5ZPBHIDaaXDteg
XDDwwUPTx9qPaKHP5+YcdQkXASRZLofT7l8w33RFEnS0Z4iA1gZI4R3fuE4Hfw0Wxmvg795b+DJh
f6UiL70C+s35Mt1jG3pOwUX0I7lr6tB2SHL7DwyxBlzV7j6g1EaVdTn92LLHR8yHO1iCPB5WqPNP
4qVEviEN2OIs08fgRWoyOgVMR5bXb2Gs4fzDd7T0+oEr+pwCdFqFn4JZOT6dGgQr0h3u70NGyY/o
xiUNzn+8KBSkxhxCzU5GrZMM74PeoT0kqQCc9XS/Z3D3xiWi/VqmHfPYHVIKSpGcqUYFfauNGS8n
KEDjZNU1qFrtFZyk8IuL04rHhjNUHhxd6IZ4GFXN0owjGzUBPufHd89uqhsGC8GLfTG8cNvzeB61
0JOE6bUQQUUXneJGT+0oZeYbdrYds1lkTkuXixqG+9nLKr7jTv9SFDqtxiJiuyNrwD5DoiQONdXX
vnU2JjJuk2tXl56LqXJGrigTuHZAg0q7tl4jebaAvZwKM4H7PABTvu6NUTUrg4bAqK2mBpcrvgKB
jLyTNaFY15OQQ6JTlN+5D5vaRXl8Vl+I/d/19zOqVknPlE9VVWJclu0EQyI3K+ERVuwhH2/sopbK
B9fflrQBRvVNMp5IyDJDqXUCdWT9DD+nUfQW5lp93tOVcQfvIcqiKH7p5+q66KkL6TQcadAzvI/H
h1GZssg24LTfCUsVz8yp7e0X3EbmEnFAUy+YfOicK7Pw2Zdj39X4IQS9uMPFzx3s83SCpvjT8I5A
w31YhKHQZYeYC0yb6/Ag68wpYZ7N30KZZ1xdmxBp9XSFOOERR4bsnQE3URdm2q4ev7mcKgBZWz5A
IITJ9uvALY8DDIJRCO1pp8XwLSR+M09GVvkeNI4U6MyCA0Z29nPZajEY89taNvyi7HhrRyoazsmi
F41tqFXEINPStYnMwwK2AeKZ2VS8AMtYw3igVUvohZspidZQ/3hoSBrmh4w0fLcJPrNjYbUS9TJ/
dbnBYsgoo7U2eUn7/xpTNQtN/uy/KRAHiUboShA0FIMHhXhEjGzDC6gKbg5DbfmPHnnkI2tHEEak
0sSkYpURyafVYaLqc3xjwKTomwOBhkT2w+8bgKiUNJOWO6+TzuLLP/YiQgEglP4N8Gtfo70mZeLG
U+Hcouy2VOp7sUTyEOw1odzVOox+7HpeP85RNi9wLKKc1UhYVOR9MBsGNfVQttUoAWKaUaRuJUxH
sUiqm+cDSqQ40wxRGc8UOHumIGQtQqISJAr2wFB8WEFJ1jndpcANkAMvH1WxnC6blYVmpvysV1NX
wqrJanqhggClT965mQzVn6av8XrnI/sB6Y5F5YdxeQQ6VyDt+nlVLpriM3daFa8BZ4MNSLWOplPR
NRySexfZ+9R7AjV7NcauPy3VcGvbGHqH/X/b/f2nC+4t/B8hVN6lfr6w0p1WOO59VzwZGcPEHe7C
tNdX5deTW3Z/r+l4bwEnvVCfZQVeuphZAP7brOqlUahDv9KQmOHGeASOkM51cKKrLh+4ttQwXOV3
JvEDKJcG/3xGUlkjKSVzdBMgjYhuFqJ9pRXuMES+KZ/1ge09AcCo9jtzR7Esgj4Unam4n8ojrYb5
0fL8revZX9ZAzQuIQpQNEICpFGeFklD2n42JYfpuwbXVtir9SD4WLfSAWG0bHBw0miXsOgs2xEaB
WUS2NvVmymGVsk9UnHsfFutWw1wN6p4V1Z6E+xrPzZlaP/ISjQhCutCiJLR+bux+anWeHsCxpNXA
0+hI630ulRk5gEAaEeECBqN0iNfToEiFhNvzGPsFy1S8rH+2gO3SCqOC65+PIrB2thgUlskk0IYO
uLDCgobMJUzDvL223GuylGQ1Lw33y47R6LWVbUI5jp1GmSh39rg/dl7NIqjKcMpLwg3ahWP8PLMo
MN+vot8iuZYNJTanNpIZ97xAsDZsbZMs9KuU4a76N1K217fUAAZYTwl6lWZUdAYevjQ7A3CbDxlo
9pxbm17l+SSgotkmlxMVNOOXSwDBkdm22VVFKw3yN4b9Jj8k+UIy26nP2psmo44vLr/oe+yt7kUY
5nc7P1MM4zNO1sIEV8fabbNdAht+jM/lZ+PxfLViBiXketj3DJhm4aShti2riHYW27XOR7IE6TKd
57yNJoyxk/yVu6Xm0MxVWdemBuMutGuLI88FCb4rdEzd19RnkNYLbYUgCdNd96n2DztXVCO9P2OV
yYFgp/tqRIEXPGfmgqR2RIut/hQ67+oYVFecEBgqOXFt+nW4zegTodTMpFMvUBcln9FHfQAJYub7
hesRmFeoSv6Z1/19BX6F1AwJxBLnaD/0Nkl5iBSNwyK5rROLYuRp3nOt+QsFbj6bYR1pRJWtuuDE
KRY8E9ARETZoTpwD+5qukbgbZlsodg2rthrCIrvn3HpK+XAon9dDz/8AznpeEghntFhOBsIthxj3
7yjZ371xBYjO+2Cr49tUf6J0PkWlfjMp+k+f4Qj/ANY3mhY8o1sV50tz/ZGxgqGMKCNW7aK34ozJ
UMuiO5yPOGiOXDLX+3Sd8COBCEbU2XkXFP7zJBnS8TN3eJjNWCvM8Uc4NYoo/WFVJ8ioY1W+P/l8
qruUKrBx1rBYiTqStSzJuQrVOtC1ADUQ8yMPOzPN3qEYlQP8Bu6T8elzS+3IqEgHse4T5yv0R18F
eYrmI90VQRWgJbvljjETdYKE93NTkhUttlX3fAFmFw3n6gK904TOFjUczhvbYu6XgHf1q1RfeZFv
R+lIUgKN6CMY0jfOiZfEO3d20xXfCPNmP+N/VviLw+oImjV2WW5LGCli759DWkkT3CYCmNb34t1D
ZMjKV+J4LBP01wO7rEpANTJWsg/xxiprVpHiFn7iwYDo9uI2ukXwv9pspvyraJHbu50nZMlLT0iX
kctIOMHMiv9/wJ2DLH6E/lIzQlVMMevMDbU4mWRguiblJo1qS917tld9q2qrxTzXL4XS/GucSeZ7
iaGeOZ1QkyVZKop6NefBrU3hT4mzoTfuA9pWS8ppKp9hv8+s/SQPfkMUR+70tp9maSHHqsGJVZsX
ltolayYED2rxWfH2VlZvBmly9voG5eSvkvwWeimH74K4SuehztgdU5kTwvpVhnMZX0ZNPApLPpbp
taY4dPQIo9E2ODFmgp1AdWUdgEIL/oJLllK5kX4ym7y+UNR+jbwWToxjnRwpTHvzlJdpgzu0LZWV
haFDOjlNmCZCmSWhqHva+R/GvGBp1pdkIspv9aoT9kFkdGVgt+jLdTtRqP0UEmBf5bAD4M+o/zkE
1GAh/Sa+rZn0vwxlo/iME+FruLOg0Lgx7CVPdFpBDWHoLpSPtsY+ybV4KeKs5gufafnmTrryK+Mh
2N5oynm6xMPq8RJUd2uTTxG8rbcv8agIpUIrcUyetodqMLnM3NH+Lu0MKue41Fj569Lb3BLp/Jt/
eZiaHydY/fBKP6b6h9a4QOPkjLVECiLESAEHf+RuAtlU4EztygnBwMJh4YLb1rvrhidaRG/b3XzG
GaWh0H0cbfQ1B+vd5Inw3T+ktyYaoz6jZsXIMgmNOVCQ9y1UHPtbNSgUs24bNS2uyKr29vYSYA7v
aLQxUZ2mQtPkDNEgjMF95RL990iRufOLbc04fZTuxuuCrSq3HL4QjRp5Bqt7dPvas7bNNBSZBiqO
UhRrCbfaFvE8IH/gG8CVRLMT0aYPEjRhOszH9AD6fOU1ZWuPxvdnHpklJjZyKOVcbLKbk/SlsEPn
z7AnTG7oG8nxzdIiWRTNSWD7QViXJp9sz1wTkai6Tj+hGguISX64EkvDDZdLC3Z2oEJsAI1MkvHM
91XrQPeMakujg4+PMYhyszEqJglzySvV1zXPgGJQ1Q2w/sIHlNfKXtOwdY7KflwQL2Qu1qMsJxYT
iu3Nilsq6UsXnOT2ipa5wGfKUiB/gjKL4yFi2EEg6kcAjxwl2ViWoojESusCYb5KcsFBkdBIp9kw
HxEIKSh1UQTbkxh2rUmdFrV4wQTHk6H5an8enZmb+pVV/fatsOdS9h0LiYxA/9w0RZjLQTXnIxsF
9kFUHJC0LC+2v01vQtua/XEEtYlajzbkSeqAeQygSuZAsGK06wuh5bC/rDMqf9uYg4NQ6oh6tcck
NkhcbkCC+1A4amYkiNtvWx6EthEAJGdC/J8jjwzYZWPtIyxZEyAQ6IbqolLhKt/bZT3dpgxSem3m
bNzeQv2JOD6hhhTiSQvP04G8dCvI/oGQJQ+mfzMWdMMh6ORZGHQC0RPsbQTmHC8CFdSDTB6jhj+x
LXcqo5Nsth/wZKJ1lJM3bm28IWo1y9kwo6MgL589mThj3qYaj2ZUONybCslZYPMn5fDosuxq6svO
iP6FL+jvh/Ec7KsX6ayFz8ieSn8YM9LaQKrjKG/HeYaAG7wQLXp7c8xPnlK29ABug4LVjISHq9sX
XLoB9+orHx8il5FBxGS15D32b4l2ELmzOIB65RAHiJvTXOpHLaowEbCaAwm5V0aELzfRl6dqWFXI
eK7JAkg5/cAmwZ3NA4nXR+iZVxtbQxMowCbXzo8OliGz6FZ8YTxcisTWKshFdnpZA9SS4xznw9MO
v+hIKZWeCoZJxxyvFuq2Ma5oIoPx0yRJW5Zep9BIbJcRZ7QNFHQplPNADC7wQET5jpcCLQgnPhYb
vDsSySVYorlG2JLAVLRrmoZ6Sluzo+QFUSV/nAUYr4+AQkUADkw/bTEJHdKDx5RoCgEISnXDUoJH
0p+ExAiR4RsYO9ffesmVEhtqfa+KPWmn8+thQUAswZ//B1dQQoDfl+zBpBUveY7bqgg+MdQqbzQR
OGgHkTeeXU8p/SoYZhSXRlLEG3uO0V6fn5tGjKNzIWd6/b0MmDQjjvNXs1Bd8ZWyAcCfXfV2FUBo
m6YDn4wENHCwxlE9xUTW72pavvJr0xN2adjSha+pWcvsjo9sg1jhiMiyILwbXDMeqrRpSQeQxVnK
zt0/B0AZbVF5FlxbEo+Nhb4tjguymaM5OdAKFKTvy8nhGe5EUxVDDtA0NvP0oyV7q4ta8HrLdoWl
OickgchKvzDIWXDKJDNW3JmNXWErApBeUuXsPEWp/cZkZ6TjglGy5YOSKc19GXG1auGdFVT31CTs
C+Y/cC2MWban/FL62RzbDymPh8CkeapkU8ROWrMKkwnIeVs9094f43zjStfBS/uC8hIs5mOnznZW
suoOiZDAdf1KAyzkfF9FOI06XwrAxaAFYIhZUtxRF9JkSkTkL10dDbmwC+mHYRGSNZ63yRlL39LX
cD57FNdM0TibN/HTCo80cY4gw3OUmqfcDmtaNKn7vANSBWCD3v2JKQ7BGbNb466f3JaKN39HoSd3
zc/ZhhNhciq7I48LyelQj/Yol1oXdrSkVU6W/V+x0phQ7kN604p24rcCKFYm3SVBYnQKkuJOwzdU
kzkf/WDM8k6dtyD7hpIBLcjqY6zdK1ImXFf6ZuoyatdvkJ+eNO7/7cHvd/jOR9UYXx4Xc91vDTk4
NElypZRPZz5fwjYyPPU32yZIufq3zAFzNLh1dRQDhNabt/Y/xNm3Au5BwcD0hGLGUISyPRXuUR+g
8eQ5+H8GxTRQN7vGYmHYLlIzr/eCMctYcK4euwZoissnuMMD7scuwGwNnCxMk57iBdBPZvkGCK7g
xS8CBAkjbbxtF03nYuwz9YRk5q7Dy0eRjUq4HD051NsQfrgiZpafZGKxuABAxoOYjfe2PmbpPfQj
m/98LeGRK+eNBj1ZALpWup52yxDU6ols/5wcg2TflN3dKFXE80gkdvaqTMIiuLW9cLMwh0fWx1KB
1VXX8t04elyff02AfGsFBBvfqLJbDhVGXp6/TO4XA+qBXl56iKhm2KY6t1C6sWtKZRiNt2+EE+rC
kNRv+gMj5SaCb4GwPlhF2S1M5NJkPoURynfXXTSa5rZlWjLhLQm/tvGpuB2Dz3ykShLdLLplwx1B
myPy2W2DZwz0tpWh06I7vcK63GDQsoxlBGhIrQeE3oldBOYyRiw67L7w7e+d9UUu9U+8rq5GN2y7
xOV+oe0QY+SHLipHOw3Xrq4OKmcE7DKEcQ+yV97khzs5Rgn+F/3l7WFrwyx0MdEBjXfEfnt05RK8
T8R52W6SD+ObfYXZ7q8n/ST0Vl4iu5KzEPbSQBw/udfbWMuiPDuqjUIFPH1Ud3fInDlBCzgWTlqr
tiesoVb/TkTZoEt9gjBbVeFrs3COfXmuUBINVDyzgRMozTTUGu95t3szd4OkagSNqpwDiCpkAr35
0tbZYFvxmCnjo8xOjEIcYziSiDcs55Kn1pHeyVf9ob2jKhdTlruSCWrxAA5zM9ACqinQvtQqepBJ
xoNJm/7tACjb9ub+i/qY2mOjxO4mAvxx1GCIRRS4Arx1C6eLLRjJrpcy7sy3Pg8mtO8mJoVliIBY
y3jLSHijKLynYX4EfjhQw+vkRe+5mkrx0kUZnGYaGG7gGo1MpGNiMUJf3pcolBM4ytzgNKLaEpEG
6j7SzxM8VB+Jn3Gv7zc8o2GWp7HQrHKYxGcGgCw6WlTybkaUF0KellJlESpY6+2pCQaHIoaNg+Wv
/oHsktWMLIzBiOahawc7Wd14M7OkmGz0jCtn6cQkVTHEFGmrV/i00/EMCGhpPPcPOzOgdOUZCR+s
x5ieV2FmQC+3mGR00bl3bZ5oyJ/74T1s960pc3VANXOGpPIfyc3zfFyfyuhiJk+UYcEcFmf+Nf/Y
+5ZuUR0Zqib880hsWVYhuNTvdKgZ9661uZZtAoVDH92ouA3lHo6JF8pdJjl1rtmrSC+4CaYljjIr
3jrjugHDuadhI2dt7B+JsRsu+0G7iMiixktjwPmj/IWaOmfDGaJTY6nEuEBnB4ImuY6o3RvUSYYi
QcpsA58qrNs+db3MiYVGERvBqlgSNvVAgrfr2JYPqdOnAPPmSslrAeZw2sqtORTzLJZJAbkPXeDf
A9wjfb0Hy/dOHURYUiDdzbl1/RH+kbAk79L1p2CD4jj/w/Nl8HY0VNCHA7oRlNopfl0b4UjwMqB8
OF3O/du1lgXBdxCeXNRTjFDJCqRBAfAUpZDSfAF3jXDGI7KuwB3LDskBUrng3GyVtqYcTkzontAy
VS1CIi0vSVB6SIj4U/3ilPvaH3Pg+2U8fPt05dMZ+7rjEEhTwJM0Xb2QO3CmKttnwwP25kciHcP3
78qEqYtyJIIQO4xicGEhqEzYMmBwKYTNQVaIkqGBcE48kpp77Py9NL4wmmpOB58owUXgFjiUeajT
1/GFNdqEFwttRvsBaByY4yZFWMS0ukalmOtusRpAG3rwLMEsa8UPxncKkwHbVyP8/+PxeUZS6eBF
2Uny+tSaH6JjoP7NJ2U3kLR/0kig64HYGH5U8z204TlO8Ct5VY+C3/kt3T5RcP2tHdFLcUpx7+Jb
Ojqy/C+CmHcbaKte74bN9os91i9NlqR5TNc1ZKiCBT8YsP0QveOQKut7jNA/BdEneUl2vVMg4NkE
23UI9ShYUgaVnmM4xDv5cWb1tKr8dSEi30KUKgWGBmDYs4kuHeezKQZcEc8QpWC6Al1paBnBxrqL
fV/2MFb+ldLaeQthfaugnyfpqcISDSJUrXwkSUEj0jpU0V4fp/3WP16xiNFhxD7dPas9tE4nPZBg
Zf+FTjvN+pZq6wO6CaU+796vIKIfqWZ7wTj7MMZUjq5kesLBnTIEKQxWpG/d9FYesZ9gwvNxz3Kg
W8qndocgU6pWci3eBrNlLanqY+eT9KDP7IbGNaS16gFvG7A5aahcomzTGMNc/Mee8w+dLkpDZyhi
pRPq0bjg9voBrTplgGwOm6Vo2qvMylqkoLYs881BMWydyqnI0Qr63cjqc8/WJWIoJXIRMDjNRQDD
trw8MBRuaWgA+4KL9AzOmtlIMHd3Ht0r/5z/+lfYMVSqr+8mgR+tdgQ7mQVPykJCkuc4vU0ni8Ze
kJyDJjQRKZYs27J/II7DFMP6YaOjfVJ9VGO9sHq4hM+EJueNJsRg+9sHV/8GL3jCB02o7SMS9t5C
h29HgT5ujGovMLq7GyCRqrhujghRiaJtJE2fgA6zl910kQpzwRi+G7TMMxRu4JStnWFrs16Qubig
E9BFhcCCoEnaaMbfnY9W54czpGSEU9T7NTQrfW8TxazKk585CYttBWP19csRfbwevzRPKX3CiLNS
wCSMSNnDSMSrI/3az+HpLog6YzIQQIAZt4Lp3DbfBwpd3lZBefOdhfTtHGey23GzAEJTeDYtlIup
BmQbAwVdbdE1xJmHdHWJquN9YgTwtnt2dypXrFEILhePltbJIbhWP62lcfv3HiFh+Y5jm4k0h3d/
Q3Vza0/aqR7E2GqLC1bhYNJvHOuVxu45BTVzY0eI938SR1p7qsxXnEv7H/0tPpdImoelcDAQUmE6
VIXd/7Ct2d7DLOCpgyfQ+b4Bq8jIpRGfj1jgCdHhQ6lxAB2kWMLqI8MLzTyCNEVStUHikDk5+cSG
U1H0v1QWlA8ePTfFgKagJR6P8K7OL3/OhBxTwLHZeWvz6AkzyKd0a39BfdiVKNb4e78PQkPhKXtE
tAPQ1pVo2SE6WBIKjNhNpqgartTEGk6z+Q5vgFhYTUJC6ypMAc0XP5Gk1JA3PdHSlylJ6GLQDegp
pVSipbfUiAnwsBAhPQjqa+Ef/ht0VSZVmCYpA68MWQeTSi+GrKenM8G9JmpxAI49aMpkVJ6P1vF9
6TnoHjl+uDvw/Pu2T9mXgVgsmWArOkVYD/KOcYYLe/8HXxwG04acarpYUYL1yqHcKiEGqaD+IB8R
v041z4/JZN6Eb1wxJ3UkQKRti0J1fjXFyiR4KHHdyj4bPidFOr0afdzJZW5xJ/olJuMmUHlIcwpn
FzD/gESBsAGVRtRFRemX+9h52jWWO/Ias/3n9ZwRNXjJxCQ+/1X3yRktlCkHL9mi+z5fWZFl64C2
I16vaaGdj5talBu71nSebgvibmcq+QWGsAeMqC1mwfE8gAFVedaGhJ1Qz0C4MrX7DHBp39IzIJqP
1CVtNiwO5jj5sMaPluVHEKwHAUR7FVZWIuK5BqxhglZSgfQaTZ3o7wEgsaKLN8J3usB9auueQ6Xk
2hUjhFOGB7FZGfpy43KCQFxUMD51BEhb1xFOAS8eI26csXHvgasyz/IG+vlf4GCurBYKUJ4WMNS8
1e/iF+myfFEJBVneDmIgxp7B1GXZcS1jkZjPhqWxNQgR6vtpoX4dDAeFRJP2pFPKImo2o7lZTxkU
+e8vbVni2iUCHgRlEfEiegonUL42yw6x67TIZHtyNW0ElJlBqP9lP36pA9u00uVsVN5/8Tx4DcTd
wYBBJDZRdYkJnz0wnbZ+bvcmNlYcTAVf4WHeu6GKbwgH6VLDWBiQaiYdFhgLfWZo6MVBzl81iG+b
zVHWS2NFhY2+MjF9JaDVOopbMvliA2P7IhzNm2gptdOGq8mw8++h9g0IzXgeaRka/g7sIJMckVrB
6yK1H3DzJ3hI2lArEkSLEP6il9RGxdqoWw+cowXn7ajR+mRUhTELdCCNnbvs2pCusxQPHC9RGPs9
FCMLYQd23Ivo7UhjokJjXg5+mIY+V86rKLhqlAL33XjyU5S7OUMW0XhwxiQsrCSgq0WeYYmoD470
lZzR7px7xIduAT/dm2iNiKZ8qGhtq8nVUi6P+H2BCa6vit9zrNJ78CqvNEgtV6c0UZDF2sZWrWnm
FFMwKY3MSdKF5QUC+T7feneIaSr/+Ot7cj70NbXCsCTvPuFCKvqWGKAn9pqW8Yj74xkSpCaNjV4P
x4M3zief+2V2fk7te5F8JEdYZ4HoESG4YoD40GqN1nCDyBIhgJBngCUIRSvQ9ofxvGaLhDLX3YMn
QTiSzt/NC1GjmWzpmdwyCYqXI1D9QrGlsM+87Z8QZUzt1QwMrJWOeujtzTYFiUTQ7qBMR/TbnMGq
mOagJy0paaQlLf2U6vhBHvEFj+18MGcbjKW3+u8I5dfUGTPY7EQZYbyMuxKZq5DDbpKQAHIh7Aic
cTewKmbzZfJWFjsenzcq7deOqlScR29W+MOOS9e/bEnsL/iRTDgTqKqfT0BDq4d6JJEzOfDayO5f
JXcTG2Yq5k/VTdLX3vXBzRlgAlbd7xl9GjLCSQrJ5ZyZY4svHJPLTLd93i3CcoQt+sByjT8Hq3Au
XIxusVzUj2xNt8HZb9UIwwG94c2TPqMBFVIFR/HV2tguNmYyJQaZl4B8j3o73xjMVi4tLB66EBIA
bCVDoLlytjjnQLupkb09sSm50zxaEVW4Ywujr7Lg6rSVpSa7vk1xz+jl8QCDZUV0Xpu/lhW6JmE7
SlnJLAL/6LaoYwZDcLAw12HCSuOeHge0H7F0NBwvmtUOU3RW6U8Qow9tqJA2q5jRCFnJyMSTm33+
7v8NUUVS4It0Nk1A2cOKXp59tNsYKLlmSomrFOeqhcdS5iaQiLyNtoB7sxA+HutbSBb0rQ+8tO+/
fvdP2FnE2l+FYNMCUlKxi/wOwow0i2RO9NwLjqNUXJr7pxCo0+z9Q60vyGxz0j7YOmBJimLi2Ljv
SJWm+dBSTG8Ixq97kqgAuE/uNuInECyfKM+l4RjQZncGAdmcnOmNCvLlcfABWkDWBK4K0x1/+JPH
mj9sm7qxAWHvhUSrqaxAdgtZOFJbNaKRaoB4KEf7hjSZCN8PoWA/Y17OtgfFlpgNZLulOnahMzZV
UMpgzFW/1al5B8NPN0YLS/Ja7y80kHYe/wfup/ZHkxt5NuELXmYsXXE3Tfy1aH6qb6s+m3vzF7R8
LGyGMY4m4sWxOLvfXn5YzGn5WyMk5VjPc3g645wGEre3y0RIsMvpO6sZHBPi4KM3hh5p/zDEM2WI
C3KVcQMw91yD2dlvZhXAHQBgbGIqp+/wGl6XKcW8Jq7ujWOfDDYlfpBHJK8F0JXAiMhh9HUk4Ap9
kZEhuyy52GHYALbO+vfvrDX7fu5xx2qA0NtEBJ6OsYeHy4HsDXiz+Hzvx7s8WgyLgBBWsgsXjBuO
0noVobVyTGAFfUyXEJN/e8FxkpK1UBIp4gTuNyLhDjvZpWwsYfpp7ZYhr9rqnMKMItlm7POqVJKt
DQPa7cek015wRoIw067IqF4ObfLixdAvHjksyvA5BcQsUYM3Z2S07nMw4nq1bfBuJ04lutf2R+Rc
+OlvlYN09dwPHb8TZNRAwtenwOpYEwqS1VTK9xYRCRqAfV7AdZtiSIrUIB5I0IRrnb97znKeC+1j
7KG4X332dldKdljEyCiiXwxUYmUNM2fBgq8Lq5J6trE04bOr0LFOgXYw3qiJxdX38bXyabuAzhnE
6w7ojMcqRBXHUvRrW6KbOmP03DV70G6vgVnhWI3dfOsCw4rcQrXzMA8I6jaSgVKxaKiCE4Mt1et2
Wr5VApwWqRn2oX1VzFAWqGXJNTh0GxUujDMjdu3esaRmcVkNyb/0eYcGTskeqjfKffIhe/+aviZy
RIrcIh6ivXFNmJWYkRTD3IKa+KeaHR2UOiInmWeBNJA/cVNaJ5zXu2y6Jc0KfSBfiknk5Z99fGy8
JbM/dSrn9N3s18lpJGZ8R+fSRc7QZVA3ammubk0A88Z3bXPw1Vs7TAyyxsaX3AZq7+uyuqB5yeSI
FcGVbU97TPl48LbjCrAb2Q3iJxdH8g+wlvj/5UxUWyOb/MMrdgWccVS+vvM1VbeEyLNn3IccgDHd
cExc//qnqQutrHyQ6nURimtqxnX2/OOJ1B+WCK74Xo9JZb8yvwkYNs/yxgnZoXld8JSwudvubRPb
n6zff4BSNVFXej7hySDUTzwx+Gg9CLySuvI3/Q+bORsni8tt3VsIGplTq7BSsS2f3SDwrS1z4ToY
bl5P+IfImYybWjSSU+qE2nt7TI9XlzIgLPuapySahOiqt09PKFxjzwcgSZqs8+6NPUslkcT2GCFT
9Jp2jNEyeeuqAZO0xOtzISvdgjTOaP4atvn+acbhk4x20y1PljSlmaq1hwEZdVUYBo46Euinfiss
f9TlUsaVk+toAsZ+kpoYtn3Jr2G5J3KdZiLte47Abr2CPxJSPLk+oaQaSq+YZxtAxOtW6RQcDlVJ
1WEmkgFZTw/Rbxdg/pWkCVUMpuJ1U2DTxoMn4lrkfPf+Ifl8XBJT3Fmhm5MIvpnmzgaoibo+S4p0
bxiv5ig4xFgRg8t+imuTt+GrAV9mMayFwj6ffMo4Hb4ntWe7dOI86FkChyyerF/AWtJGXlxy0UJQ
w9QakY3g84qAiFx9+JDmj5Zg5GDdxyzNzJWguJLAb78AFRCVcufO/jSE6FjJMJ/bW+QMxjLgPr/P
ed5IBgyzLaH8yV5jCZv9PB96XWsSYr/HJzqUUq74aw6Kcsp7q1FLeUIEYAfo2uk1RrCSzo2p6P63
ax5YkGuKUP82CYfMb9lrnEIutFraKKJ6Sy8UrCVBt1I0W16/sslPFqDhsZ+0la/Fj7xQFH74Rp6a
aiKDrkGdqh913oExJeAzpqGZG74f5XrkuXr8TrSTmwk1LJhJmnd+h74WeuIEq43yTy9m6Gv7CNMZ
cHQf445gI+DX/OyLTxpeN+elwIeR3yG0LuAHuLu/wcns2AP57FT0Qqfvx/xj/F56shyOIIx4PTYE
ZWx5OjvuYkkE41/q63LSvETIjmqEJWbs0FNRjOZVaG0SMpv55P/vSvTQaWJg0G9rE5MANj77Wbw4
AhDxgAWIRYZhW9FfHvxvfH6TDOHvZM+6R8s2ANTr8g2dNFxcl3dyjJN+wz1GFvkyxT9EXe7Gaoif
Hul+K75Mjnz9Di2s9ry7rNnnGHZ/k7PoBcI0olF1o8cqr1IZD5zPhUhalXwNs50tskkJiYfN7XdY
i+DqguzSqpkQ5ReoZLAV0mj4C+v9hi9+5xknuXf/6sf2/BXyAwcoACMFrxdKnAKN3YUpbX7zOc+J
2cOOLbLBMorohmSKiUWmjwStNaIYhy9XLUyYNPc/+ffQsgM/7BxF65bK1N7sd4VN1H2q3Maa4kUK
46qDh/LnHnC2A+CaI+ek0opES4V3Hs34PK+RkXklKY0m+TYxUPjQ+xHnBpUVoGRd816S3UQVuBnI
QOg48ut3jCHerBo5Z/9fgDhCK/njxOz6Q5PigEUUXqBhPRiw0OQN922pZh6XOwoUuuWwJuu9tf57
l0ZPeRzoQw7BT/ds9G7Yqr74QFQJtkQeGgzhIzXouOwz6bcX7mv4ZYFsT2ljLT0oNsZDmGWIoMGH
lGt49EOXa1ntHiEANRtlBZjsEVio1xnAgl38kxb3ftqH6Iujnp2n9SjqtQEa88q466LLcLg5i/Vf
AXKSX40zCJzMEpgsnniec2aYxY+7Tx8QKm5D4hkm9T8vYQyp+aekNydHoUTdXlkywMrOpMX+eubI
9Erl9nCxlKra285jtkjWy7xKRHLJ72FPdPRQ30YlWoZXIdlWcbsRgw28zGF5R54sxSTN4N9J9HQa
KnBfEFCW1DQEORcwKZ8zFkzf9dqYXlfWjRsia+Mz3pZF+P9jqISagdaTVSID+9bj7Kn5mLbOsHna
L1eBJaj0ciiPcbh/01gUr2gz2Ear8jG28l0EARWEn6Ui38/jDETd5mxCbUCz5RDrCGcNQtIcQpkY
NRKJC6NMRJcR6+xc3aPhAA4uvuHR2FEtPNIrnX+snmIvgCGYDvCTaRV0So0/JzYv9v/YdCGSwVEi
jLQ1OWSl4w0PnSo29ny60mpLeOwfB5SKMidC2KMHS2blIe5qXfVG3WXh6Um1/38xjZFv4ZT07ytj
vUi9YOuPIWE3nQShrs5f8usShaHD2i4c093otCmVMvQzeYM7Vfz2V+XInX1exAafWCvNQJ/TvAW2
qyR2EGo0FG+RKs2QXHF5ZYzhSjMU4/lUqwveBQVrsW+RUYmtwuvmU01kfmEv7GQ/Rd3G49QSoJvz
ErbYpT4zdvpUUl67fdIXdGoSYqhjWGabWPFApZ9zi/etD/gbh9O3ZUeKOjXu2G8vLuVL6/yAHL3r
i6+X9NjbBlDJQMvi69ARvr8Vz+K9DV5/rhgfICwdY0VcelbWr0/EwbTNdXsxZ7GMQaa3a+RaGmbD
Sj8hbj5AJsZ3hMiQzuAFYdohxCZze5OghiVIdLHlI7siAtxtK2Zld9uZsdAq3TFjVtGxYt6JZ1Sw
2DBjzPkdgqKZhlPTgGyDqjTcWKQ3JuNbgaDvD4x741PaqczM4/dE6MSj9n30Bzve9cH7qBQPgIl1
KGUXDGlvji8CVgR97u1zh7rxLnClQyiUS0VPJXFnBqOAYbOYmx9zPP6HNw25T2RMmOZaxzU/hDLh
3jPMHzpIyqZ2ksehpjN4SHvFGsSMDU5D+H1/0PYTG/zfmsfByAvv5sbN1rrqWHI038KqDz5yEhmn
py24krqg/ui045U2sSwmHd3zyaA6WoRnEuq+itQEUeAzWdYEt6et1RnwahkmZbhASK0YBxV69t+m
BJHOn7UYTvJckPJq/iZCBVhSdMzhEj8+5bRof1UlYPUdXp2ptbqXWS6LuuS6rNAXkeu5CNEafVqv
DIYDSJeRsXpmr+vvv8rlBj6Nmugebfl62dQqN3qK1qjm7pfdtVyR9zh4Tr3xNwFBpdZWOkkdXkJS
4I2AXiH6yTARhHV6gYfPkzmBXl/Ij10rMd/tXQC6x/PsMPU02I30xAAs7zPjPPYu6gXz5snOUFL9
gCJ9vaDVw4SBabERckvOFrakSxBLJdUhvi+b3WWEYcQcdJiQ38fc/iwDFTQ2VZWV6Q7XcbfYuzuF
Uz+asavmXoCP77HUiSuLITbI3bxg6zz+GHR/bC2C4znH3RV2iEzXDhwjeBKIy8U9uyF425vfrh5m
LcKulMlbq5uAwSqMy4VVEMmaILrKLF7bSnJR2UCGI320hJ/mLIjQj2zI0HhYnVXL8rbxj0VGGZCc
x0F8BkovekbXPiBZbVfNaudP9ROZMpxPtjos2vjGUWMIttiXb0PGT4CYqP1sLhXe3Rt3mz0Dd2M6
NUfpNTbdOl+oTYoQ+AUf7xdKfBExBgZ+kb9c2iNUTrE8TiA+GkkBb129UuLX+OxN+LLlSfphlKlA
9x/DsAVwUIwk8qPvE8W8b2LIIIwuq+zpdF84MzHNz8zFCAZ2OH8PEv5kqMGTNWI5rokR1hnkqBHa
Tvhik4UZc5AO6AsFWmKecwMIA0N3P4XGjdw0BB/n3t8jU4xoGiCscEe2J8P8zvk5bY6USUq9FZKR
P8txIFDhjjXdkevt3Dh/YbFR6W2lPM990nkXIPt+VL4A1acwH38Zjl/yc28fBbMEHF+pfve+mVi2
KBUbdGiSO+6bV43j8wlMpOq/J980HjCAQWMsJOPiQBh+BO6CM+slL15xmiPqqCCEvsytkP8syi7R
88feWUAFfYjLcNQWU9sf2KDVpG/2Kev8Coq0ADjqUuHg3GoGvvzG+pMnta9kzf3CWDufJO89D6Xd
gZ4FfhNNT3rJiMBKx98dmPgaSoeIfqYuFJcL+1N61bGyKTgxhC/DdWIRn7XFD/tr3Wll8wtF1rUF
+hHW5HACY52GYuB9vnA147aQTidczjRDSUM8+psydnASJrIzBloGjNLxOKpE5hj/taDriOpr1Ymq
cz42EySGoC1rFSB6+EuZxze6Ukk/TceOadNrEzipMdkW2cdCF/7CwR6qGaU0wKOUR77UfA5Jd7IK
mrZXAp3cyNCBTIx4klDJZRLNC9bZXpz/JAvwoWpzc41FimZ/osyUyOG+9eZPOq47XAbvhR71lEJP
c7hwSnzlYvb9tdnOISzG6W7Ip0pD+m89/UhA9c9bFhUjFCSjdGy/NN89AIq7GeMGIVrJBQEiebvl
T10jXtVcTHlS9pc7e87UELdOa43J3tfSnt6iBFF/eXY2YuQo84iP9RHL7q7tXquXAWPK++n8wKIv
4jU6eq3LdHI6dT9kVbngTC/gF8AVIOLSzdqDfYmJqnsdC6oSINoMrXA7mxxSSRuYXb1lBsaE2/0Y
e94uV9qL1zEyYMmhmU7/2Ed28uwXtd/KA1J6Hbhge7ldk0EJnbxr4w8yOBuOl/kZMbR1UptOnGRf
hoqaAVUZyN6cdjc7A46aKgYqJywhrK3KdbOOzY8vxjbx309c6OnvoSO/lllzcTt7E6/XzaIuGnEu
oGOMJKelcPxgHXjUO7uqq15xTUcTLPUYGIK8JdhVb8xPS9iY4Z++xxl/2e4LEfQo7FibQFrLPYVk
GWoeL+3AoIsQ03aQ8sh2t0mVX6FWRjSPcG3t/j5y2XOAFcGfR00srzpF7W+GrMvbMEYR6mi81pJC
FutZFkbSKK4ug4UhxNN+3kKD6/oYJhfFkKFREew6GK3K6GPQ5ck970y0lb7HknOZirHlC9fpTnGS
wTwVUBMHYml95oKyhu9VZEmDUI44MGu+xkl9R9rEyh5P6FlTH3VrlhbB3aVbBCaYYlLK54sLKjO4
WfgjBUJvtL12BzsZsoLzj/yEZHhemVk47H2hG+EpZC8oSx3Czg/eoz92xGWKIydAhjO4nV8q630f
aUd7cAWRDZ9lq/wCpyGt7UbvzwPssPwkYocema5nvg3szhPNDKnUQW7m+aG4c+9pxjXgPXM4SBLg
ur0e7lnVFZJzgqyUdNVtAuue+DMdGI6VkPrv9R/mrEYm7upILr6I0cvdmYggF5BCHJ/lH91OZ0kj
hRg17KSZ2FIKC0ygWDARAo3Rr5JlKirNNChi9yQuXgTD/3M9eUYjeJiYZhO4CtIajV4bLUi/nKGw
QvAimP9tFwL490ezvDv0/uuJCNAdt2UTkMVtm4n2E9DW6QhFCAACQ0EBCe/+QECkZGvHlsd6+3Gb
XnwtKho3Rekrjws1P15bREPBPNsdQ1oOu1TB4m+KUJQZJU82sbzmP9W2U1GWRdPJw47vnR6C01VX
BSyKfO606tGnBlH/kUAEqkBSry1Y8+wNUd0ap/3RBttgb9qvosjw76kRB1/KquNsLYQNRuCXq5dh
v4InE6OUU+CfXXdojmjFNF+/+pepdY1qw5Ups4537yLQVFZNnKnJOhAhmaD5CDNguD9zkZ3NJepG
/jMeTZuJGpcB9TVZeNo7c9dCVI3oLR2iZDzJatZQPmRVFcte9my12OJBvU3exHx7XbaOm+NNcDN9
cszB5Jc03+nLpp9BPVk3g7TxSdDzkU6OIsAm8S7HLObjqotG/rhyGJ09jtv/GpS51s7JP1XoImpu
6O8hZeyXegCYmDHWyLD1/FeThTKiuyWUkgFJCq93esryrxHY6VTiD0SbBY9olN4oLKdQqj/yNktD
x9lujoneIPJzwPr5s+U2yZ+x4XEroVE53dQwboPMOE8liKIZkgkmk+uGBKTpgYvOTBKR1+jrKO7B
A9mDBhwsfkOK6ZR67EnzgMd+eqHm1+9uP/NNj3Mi/R1BRquE+gq1TsZNF4QeiOCj8pZdj4bvro5Z
H71a/1V3WXfzuybRJGhWXw75sH48yL4B2LMfxLkLAz31C0kt26P4P9eNsNXog1y9etrp6xS2ndcM
4BlpYIW9yC621aVS+UTYJ9bX3UlivrnUDysBxORC8H6QEHZkoWFl8gzhLMiualMpAJzSApb/hir8
XeQdQ5rMJefZN6FBInRCUW0iu6Z8ArjoxNmlEC7lz7lIFiDtR/woEif5qj1MKwvN/mac5VQWfAe0
8BeYiUsgeie6OoDHeanAONJ/lV+sXtxNtw12K/6pt+pWMcZFhB8thyf010t1gu+9Hr93PHO2vZjK
e5J9BeXglraDs8Vfb+jnY2jye5L/7P7oiOgLfFOkqNdpfL6Roth0mhWQGTk+Z84cNdrXzJgMxoym
UpwohT1Xu+S3ekd4OeEAbgEYlg6OzuqMh77wfVUZlxEpuNWKovhvrJOIKoAg9VyOd1g/GcdH4GIo
F3sFEiTQ4w6B0alxVjgmVrhvzzk3AQXg53blJlqQ5BwmNbRLS18JZ52MhQnIY0ng9r9At/4TyHrm
pb0GmxR6j0MavyT8dpfOKD69bsYXoDA634Sys2bWw92IHE4TEtZbDO6pAOI+Rft7pvmLxQ3beQoM
Cp2MLIGqQc5jWLtuHexaD1zdhTUY5EUzG4s+1TGGFq2twbEBssTM7jBnVFbvOokpOeMw9HIEUzpz
iWNkHbsnI9q4e+XleYic1ipMnAtIDZwxfNbGEcZXtDh7SCKIw6FnR6e5CdKHv+GyVlOQyoU/hB18
s0mCMMn5TiPXFVBP9viEDo6NeNiiRPF3NUlagjrVlh+FwFsyl6OefVq514CparsIxCqtGYZDrLN+
rI9ZYF7M7Ud85h1wFK9wQ7C+U2XzuUMyXz4h/cz2OZ+211N2YeHe4L4/59xw4LRdD/z44CT3q5m/
xk4AFRTnzHmWMIjaFvOSZib6CNKHDmA9iaZLk11QX6QS48RFDpD9Kh3xTwX+xIwX75bt1aBrgUq6
smbLRgCxiD26o4KWvj1hQnlgj/VifJgqvrzOvXYgo33sPKh1MmY+OR53cKWtIb7kfYr90Cn9jjmF
CMNd9v1w8+w5Y12iKJrtM/YIDY7QI6UCcQsqC7u9slzvrLbQAuGP30vy6htaGmlK0qrzCIobhUQt
QvpFNdrml6m6APt7o/kmoJPqhrh4Dw+zBHHygRIwpOCjgfSFPLIQxTlBZuo3R5VsUQrw8VlfZ/hU
gluWZn4Kh3EktPmA2VNquApT/CpHu23k0R0TsO+D6uGTnKaC0abTV6Sxj4/RYisRXve3iJnoDAeS
hmMXEp0m/ngXUbk5kTGVQklZ7R4W+E4mPItn5MMmnHMD4VWYimty9yS30FfWvWopEsHNVXNvWQwR
L3HPYR+6GY5lwoxIBo1Zb1pOky4KMKbhNM7a8K2dJAGx/N2+b30W3E01c36eP/whcv5E8v3HzmS+
hSkkwDuHR21a4KHEcI3MyTi1wnuee1WqK5sacbKEXqUIp23R+tGdbspOWD3D8Y7E9lagHXt0Fw1r
ruDA6s2DBqQKFBFW586PVFKcIrS+A2TjvVRxBmPk5EnqUAz+WAE9UzF1MOVI+7ehCBGYEwKDTc39
s6PczJ/npX0HhgEagv8OL73mikxpj/d9y+B22PXiHPuegK2ccwHoegyPlsrAuBaiR//ZNkFzs3UN
uKzcZvFj7Zd9ZwuweYuC+AzZxdgE6/B0sZzzLl1n3FCV1MrqV+p9nm4SAFc7DHEUiGdXVaGRPtJf
ZKDD92XdUZNG6Av5mBak2mDA7H63sRdBgy6XNxsXq4vigZ/aBJ8QD2UOs9Xj+oNp6HhZi5iIHWzk
Ea2Tg636iNXcskz4lQiNoWPizxAYHXX7eCuGSQ1jO1APm5q2669yA+DQRy5o33DLoKNSvTwLkUIt
KPYWNhFj4NIfkt8q+upr9AQocrfQs+A4U/d30HWsaSTdarq3NjYvS4BFkENros+Q8FExjh6qjqBj
0g6qIZdyCi8vvSbmi5poBA4QCDwLn1N/WM5tcu6gLR5utXkXJpK9yOC4A91nPzbJPril3Y7gDePm
zR7gvqmCJngsN8uO0LCyxwHRHhe8zfMftWbMpQiTMbqq7jBdoMZQobyl1eslZb1x5OX+NxdpEf7R
LM3yl6FbpqvBktEWBeqoXs3D3Clz9JLQoohUlYas+pD4WLxo1pa1r6vpmx+86AfU2dsgDmdk8Ltn
uhhaJceZkrs4cf3vWy0zzd96Z0s0kDb7EgMr0al6RmT0qIJkH3JsndaBWiE1XvjdnC+CeJJTFpR+
T9mlVWkK3ofJlBzBUohzlK+KnnVpGj9fW7xDmRCHzJUzuVjjgIMdWslrN25X61AWtexeNYN8mxRy
0J1blRxfAZQro8pgQ90H9Z8gDa2lUHzURFxoO/jMq20ij7SlS3cnd5LGDuUmV92gMMhUGC6NlL1z
qRNNCg/j6YpnovVJNcJHKZJZ0MyzhwqC5LrYgMr/wM1pGiC5ukdhzPkbwLF4pPA0feg1zDNxQ4c9
zM/YcQKgWcp7chaoc7yXQMQ4SVF5GM1sOduTLdN7XPJUMhx1guG1R/WSsJxLC4E98DgbFbBpk8Jb
K6JetQQ6XH6/oAREMUH4WkfomV6z214u4gzCQIn55j2wHbWmDeOBwi5nhdh83fvU4nlyKNK95MOW
ZmcoFtmd/AoPHGuJ7DZKYkBQAGqPnanCl+Ngds4qp4tULVJ/UnqEJhRojLa8Kf30nnqErBtj/fkZ
dzJdsEzbMD9e4Xel0hRrFQOFw5zbI7AJWogBpjAgCFxKEmAQYlFYR2n5w2lkh1PDyCMghe870z7O
0emtBAkHGxVyg2pzLse//A75Nz4lgUCEcZh1qNazI46clZc2w8DsRdNUhwicUnFbLUamfN5sOH9V
QOICzDIU0Maz3xSesaGhtf56GhdOwW8mnMRzOj5py4jwiiiNzN3HQr75pp+c0WD04ri2PtyVl22c
/RzFsLjOleiJXVF6ywoopPzzlzfla9ITrDTVcWcQHztNwL6mrDjZ04v6SHCHhwlHHpBl2dxwpuHI
n18Sr0m2O2YKv2loD3lOrtWM+oQpmvEifEOQoi3vxHRggy3iie/wyQoEzKSxlNf1ulT2Mq7Ua+LQ
HxBXLbJI7OqhoLuYEFu31xzm40hzKa78KcpWbzLRMTAJ4n9s7JRwoGH5Si0T9L/iHc3IN9k+M+NS
FpOLvNzHKvJWmo58kMMIOpewf3UEnvkhV5DZN1yN2s7MmR8gNER490ADuWjssLx0u6WdH6PlqjMF
hYk4rgFReB4INALd8BhmBODDF2zQhzvYxWNuSC4Go4Pdv5ZT9WR07PeFAgfr6ldz0DMd94DYWCpM
H1pfUqHGByLpDKljMwGJH9N3TgnsZZ+S2qpsxE3Fz4ulu55eTCDSIZ8Xt4im6LtC5dz0RvTtOkVq
LMljjTPnC1asuAF0r/vsudF8FFYNaVaqQBt3oQmozWJyjmEJ94XDpv6mKP0rAr2WpK/LpdHMgZen
0wb769FcDdh1DXN8H8pwRPeXimAhhcnk/bNObErUgdb37hFG3oy0q4K/civMShsmAhenufT73Jb4
PDL2Mh6hxtverYmA9NFoM1fPzGRFzr7jH2UqdObZ31SYyu9nttBx5mP2haaPAadAPkdeL90r/2NG
e1uTdo25UkkGXuji1TNvFqxrSaqnDeOtt8Sl4BV8NrdeOmNSyo+U0uf2Dj+JnqJdbHeJs0kkFPUg
Jxe7+AQ3CJpwZ4/L7APTBAM/IgMqtIEJu4ypdEvZtFWZXi/9azuRZ01q1anMIPtRYBJH6iLbdDvG
YoBAtJJs6rTyxDGWvlFGtY9Lb06/r3WeWqkclZ4mqj/Zh52FcFDD1Kwxdl6TOmhxhsg6XpdFYEo2
I3XLqg0KSAIUqDsBZTFH+K/2SrlcC/0gDK/Gx1vyD51DEOg/1bFG/kuTkzMqOoNW7HDGMeeUfOne
YCBZKA5fXn50FZrfWiEEEQJ2irUkVgQSVSoHsU7KmjlJmDJBhK5Z0DQqp3P5xQouqS66v8I2hbwF
w4A8KNM23e9c2ytstwd8LwfDGaoUgbMuG7qirTgeE1PA7qm7cwhjIGtY5QwiEGsJjC09HUj1ecic
ReMqvDnkeXoAYKPSEi4SIiuy3XqMcjtX2SZUW6zdhzkjJ7P+etYCp599l/Np0YPM0RJ/KJmoYQ9U
V+wcwsDqb8nEB9Q2YCOkjKx7yVWGC7wopajs2Td2f7PP01wAX10ZxNgmJLDtZ13ExPeA3HMTw+gZ
4SXCCOYEOh7bXZw8JLvnX97qhGzgRgiR5ksgYnAIoJBVskp0kHeRvo+y0YIN3wh/HOu+/QXWbHm8
YLZawlDZk75a26K15VIaUrpBqqxc6xJe8wFqTlU/IXmADk3HAAWMX/LwY9xFmj2C1JmlkMU/dIbS
1jZ9OK0W2UycaF7sEZzAHsVIWqA3LaB3QWCAQc+K1YIUjfJP2W2nhxFBJFz+96bUSozbzAI9UN5i
bZtDoQbNBsEEEf3ghfBECI74Xdl5vU3jUq/bizwwPaCThbs+2PGdhcy/4ejAUmk9keU28yBN4B0y
2MtXINckDSTIkY8C06LDJKTYrTFc5zA7O4iA7sH/t+JKwu7xWYUd1cF/nYe5zIAHzVlY3GdGe0Uf
nD1dbC2fwq1h8HHH8/u9J15NJAz+ZALcJvTP+KAonFX2zwzfR1PmZdQN6jeRg0SJrimxt7eJtZqa
5ve6Qh1BIzs++wiDwKw1jR7xefECmFdfQMWcSMLzDJSBiIDpuMnjnuDabvGKFvF8vW+MZs28fzb4
Z1yuFLloqJb3hHUXzOS3rX/W0UDqrH0fpDA1e2DOyFbPOTJ2+iH6t+HRXDTKRcUkDBAKjYo34hyV
VMivm6cceyv1kcKenhfV7TXI2sGJM9LpUgMfxVz29jvMlLftNWSQYffnjoV8ReogIqYjvYcLvfhi
rR5ZBkFq1yTNp3DhAneDUFB1sItIkgxq0WnFsUv73gECGS1l3aLDH0oz7DLkIL9JKZmTb9dAkbiV
9TDl7QgQK+Oq3z4z2OdV8WBRiP2+FZyyg3KdATJ5AwuVIcqBFsmUk4TFl0zH5P9X35tpku21zILt
Tc7Dw//e8axx9WuXmEeuNWGgiTES9LP/ex90qQC4HlFDgyP7pAGMvooFdjYNDoeB77IDka/HgUgj
UuWeYiixkrpulAR5GQlq9IwKuw/EcQUl2l/Cmzulz5OokQ9Dr8R64XYQ9lgvxeQzNLCqkb0ZsYNZ
rgJ6izCNN7P0Z57/Z4L9Ed/btRo75Q1Sv3GMeMKnI7Xt5KqsvgISxe3MHZNrr11EfZCTWBSO78+E
EDAYTwGaZZ/lC542nHL1ndjgI5iS0OINHTfvWQfZ0EaPmnQzKf5SLnWHGJfKxtTxCvbswqSCISJj
j1g3SgLmSMExQSv8s2IhukX0EkJvVR669qv1RTeiLjDHNGTKUxqziXEBYju3w/KrSki4EEAPvd7e
wnCiQ83e8PhbxzapbxnXd+a2Cf28ruACKRW0ljN3vIwO4r4F+IA54Eej6AKJaJIClOkfEnZux5b9
M3497P7meAp4n5c9uEu1aqxO5G3Nf1iStVAvGrtlY5sQhgjvzy7VB3Q0V0YfU4K4odsa9wudUNMh
0YgXwG40MndA4C2FvIBc9Nz8TTo96I2CsEQ+6j/6mczUWVz24WjcpWEpANka5q0GX9r6ffMzKLEj
ohMHGUarQaZI6UzwgLbHbEicb4JpY3EtLpeIw5K+iBDduXtvG8J4IAU9NoQeMhCyRvuCsmcBKxWN
kg3b1si24OiF65VtHLL5Tq2F5hmeY/oAF2LqlgjZXXEKDUSvqBQsVr6fTnfVhPDE3aD81FgxndUB
UElo8WlH7rBxUqmLk+8DiMw6DCg7WADR0XnD/+SXLFuKGHnjQh8lvrWsH9SzTzslkeJrSO+EcFbK
hmA2mnBDnORWMLOWjgxoWiSWIlQ2ue2Qlf4xIe+WkNZEf4Q3J1G0dfMS3f/yi7QfJDOrPs3M2+4U
sRZjBJ5sfkdW2Ka2D3O/tUkFFmTTL8Z5OYMHuA/UY8jHINspfIe/R1J4NrSc5SUrcLM8CdQ9uKA1
JfW9ppEgb+UzOhHY37H4bvlA+G/ItngTEj7QJ43IvaW5kTdXjTker/mkXSiycRMIcZCMNbYhS87X
2aWTGqYo1Emz11HQUZi7+4COLEnhxCaSaFEznLvFEtqyGj1jfnxvmhJu+v4ldORhMwoWaJ+kFaVa
wlP167feXidTTkOg35fVa7m9++2UKKXcV0uY0ETKmwVOdM5srW5mhA7idm5UgcSDT9bva/Y1SmlR
FaC/mr+Gd30G8JsyF8J0Q5MDwGZ8uh/jprCP27XfPIxywHmJnE8Tvn9nttJtobs2W9833cVwWYkY
QZSOOIv1IrDTaq5NSE+m/AbwVhcIrLZcsx1NdW0XKbskuso752Ts7QGQt2olLVPYP0DqGxHkrwVo
fg2dGkhiEa+nNWO0wJrGmTwdcixbJOyf5x30bhtK9Xwg/L5biKz3omblcAfULJ3RP2aXMi3hz8pU
WPiokhS223kJSpHo7JdbntcCHDFTymV2cIy+eB/ZjX1xGfLKDEP4JzAcrVYlAOYB05svyvjjcTDU
XXYNHN9TsynPK5vm8BLPzDWi0qnf8k498ckUhSwb1TmrSHpbSW7BQRTgInWOoezLRQbf+SjgWmSZ
jVxgPo5MvmL/jMv1rE4t5n8r/y30Fs0wcfT7Sf4agTdoIi6Rz/tb6ZzshtBssLvzeoLmM8C5rSph
2Kqeh/f2gDCg9lj0AzWEDOM5KssEUTz53IyZ5foNpyl/6xDAbJeFThsmgN2P3op+kDeoKeEcC3ib
oErPn4rqOS7kxrwsKARsVXIdvTwQO//mrBFqc0rMxq5rT+5YlgKbrgMeX9iqzRCcg1mFF8sPybO6
DfQo01sDFyuIwcsDSUFyZEi05FRZ3Xlt8JhCnNLI162F/ZMrb4TmEJ3QAP2qVj1zyJiKVJVDZtld
7lsnxFYW2rEo/nzP9twMF9H6w+Y4SOwO6xRAZ13rwymOmRVAIamXFpQl6yb96IoqLgf5AmehUg1Y
F48057F2LY0yPoNComjCwqRw8qD3P61hzAhD7UnhCioBxThMz2gJpgvV5im0g6QuTXP3BfG2EwKH
dvp9cqonQItAuJNpgzBAhlkglDLhpNXjbbDaxdqCPkBZoOYPjt6tk7DjO6ZYMy4mLkB+wmNOJduC
M6cmSwAihVRonbgur0plTbYgPcROKe26sSmtnuH99QWZVIq60+HRbS7rr98evOX/CUu7xNI/sPQS
k9wLY5INEgHrMzdL/1G7+5MSxR5sb0OgROLtpNNtzdkLfr9jcrjQHyb/X86ZYPOJQbtHnd7qIsP4
2TjnbgBweXywvGGIHl/Atgcl8xNNB/p4jVN0Pt53VewpCNyiv3gjXzEaoZKJe1tD2+deFHrVxADR
QIaOMKqY7VZRY6OnaOHo5U1x3Kv4TROZ8scm/SnRaXG815M/BSBVHPmccH0djIerV6P0uLENQTX/
Jm3QZsMgLdfvPrJXDTL7PxOzkyWd17RovEwC9ykUzVERYnAuhrcEklbEFu60MCrjUSgXz8GiTyVj
oj5ULZOumojD2Udkz619lPphb0gQ+nWblu86kypP+fSLtWT7xmgtT/ad/LCveq7KqKKET+c55uhb
KYE/HVjZiBqmBRs8aIWuUDN9SrD1TIC+SMdQRY27DwDztfBMOx58qwEVqZ1u82GFod0wVJJQ+7ot
Xs3shFBL90dRieV3sIYo38nwWntTGM8ixVA8FpP7nuzapJJlrWaQGaWem40vvlRpLZspjcfNKV7Z
LwugI5jlGnpPQ5vzvMNYPI2zcvZhGIYwgfiToY+o6kFY0HN3My2YPWSwRDSmYU+y3Kbr77wM2BIz
+DLfvgZ+8DyvgLjr8SJ+Nca6uKjjY+mJ/0oyqNWWscmsenox0lM2fYdzWBun6FfMvJmh9u46CeBl
kAz46UENy8taalP5TBY6bfC0ohduMsaB8ExJdaJIdTunbNYB0L1VJ93LJkCXv3KYtmliF4WgEk2H
W2lnkr5JDCQJx9o/VV2br1XACZ4kxG0g4bNlqq9T7XxmIWhht9ePwbMqSM7hUX4StlS4ZB61gs3a
vAswU1Hh1Apq8m4Vpc7pt6FXSXeIQ/B2E/I0X+RJi5kd53wxIASGsW8oV21AqSeoh591vAYdRlrY
DpQCCqXSMifFXu+sVLwbxAMRxe8HM/S9hSXEkCsTLzbSF0yzB8GYXA1mBKaAMnWBZxPnmEhetN0B
XYAUcVtuGFj/mPJ5OqXfnN2VODuyYbpLncyKqtDmhoHut4XdsSZvJ0ueWrGne7rljzx2Vv6LFUCP
yOfDI3DxSbOHWOCJOSbrAuReH0QIMDF8MT/tUMVsZOfI+Z2dI0R7PXkZfbnfOxuGcmFLnb89g1GI
w2ltZnPtv9SIQ3XuX5ksbS9yeR3rmfp9bSk2CnNtEOoJvtNPDLR8cT/6/tK8H16BlWkLLFYuL2+g
yViLMXB8XgYw0Y9zGR6lQdWMlCs9HQRCeT0kHuzkp/HKfeRgmcZp64mrDJXREWyfqjGOehtli+Qa
Ye1X7Umtn2bGa/OKNywmStEzRjqYn3ef9aUo7eBNYSYyNEWaV0bSkNujJ1BjbIx8V7v9+mbKQlEC
/UqXlhK437FXyEAK8Affy9Ia40Ox0OidURMgQH1z6UedQOPjoJGvovNUuzhKiugYqBhooFt1ink2
7AGJNo/3wR1fuAGkEkAYIIwh9kYNP/5Sj8O58kEp1aDsMw2Ep4Z72sMLqrsHVv+/vzfHGdLjImzU
+NUqvCSUEhIoVrs+4OlGWfjuBXBIGufFmkJ+V6YOt7iCY12mT4a/3akfBulHP0soKZyZr6Affqu9
OneyU4/vXfF2OW8hoLXF5GpO6N7yiPKZwx0C5R2GI0vVIJWoL23f1uMPrgO5OOXUcRj5tgRxZ7ha
VkgbmTvtHh82Q5TwrHSo7gcozvBBrbAd8CoT9x51DJSnDRGejEibWvxEGnVCYrYSy5ZXNAOUrMNs
AOS8ELD8kjtRhBcCTWEZa9xAG2VVxltRqkjfZ2Nbr6fekgb354b3OyGOAnn17UEq9P6hGC9jzTQy
iitO4YGdnRV095m8cR1koHKWcsjonR/ZZ9i9AJTHzXdjb31TCISvOjEIS0hlbzibyeI0kl/CfSGr
mUMMPk+Ot3UgcY+WvHW0Jxy6QXugvQWmhpI8b0AkateGrzlkKJixIqbnitW5DPzpnfydmptIGCiQ
unOvfMMO9SaMyQRmqY9N7G6mUgsxMfWT6AX8XCmHHKEhoaAwbEGBaRc27HT6BTky/VwtMXbcGVfv
P+xYIbnya2F/Llli/9TbNAVIVVYZqHQYjlSV37Bkj2gl5h8Dy0EU4wBw4bKOqhSh9PIt9FJUARy1
cbKTjgXkcUTOu7GoZAldJx82+yjc41e+OXz9cNuOXpwdw+Hlqm3K3wrYtcUdpl0QuDL3MJvduOD7
usl7R1EjqQ89ue5ljQJi6JHTq9qJu8iQqjs6M34Y2duT5FgoRjNTfQa7Xpgg/1yRIkEX/BQcULPt
RzCXGrxP/qHnh/fXc4wqy2C+1LXL++lxShEOCwIqvPd8Xz0211BOk1O/f6dfJ6eDR1MYRKH7F7KH
eNHNWXcMw6uCopskV2enWgV6azKF0uCbs3fufaUjlBlPUIvVghl+Ydfl5gCg+AM1VmW70dYZvu22
85MsbhoUGGyG8kKPwzX4jKuDkvAE7ncCh4FklgPOGLwHpcqQ00yYZamRxSVEfzH2N+COVNq4yr6v
gXe6ANroVizlPAYdM5cvjrAb89PFe3oofdMiMB9M2SjXiNBl+R00RDVogak5C5AlWfLTt5TKD57p
yF+6JykODtyRqjWZENTkZJDoxNLkzyeLGkPsOMjD4SlR1e2YChNUpbVTFvXJDqS5UBc5ef+5O6e1
NzdQA/xQCdwGe6FzaxKuqDGCAdRVjDMKxevwpN0i3vg7atMBIqXSimir/IMerNX0REvhdbUZtlpU
6YvSNS68SyQmTxMv3kNxc2QPn/mr+EIKVzn/3lN0eTHQ2UhA2xSS9VdxVc1shYYXt6FmMFKS2ufA
siqd5ppJlCjZg5KP8CgovKP6y1KSDJRDTWBo6sMHYlaxzI5EB24kY7+u00cHQIie3F/jnSUOvJ+u
B9VoI2gmc+3KjqWJcmQCdsJ/9+gSq1hxKagMglnQnT0dX85Ckb13Vs1ZOYWiCC0sQmYYyGdqKgo5
VmMwQkiYy9ePfXdZDslBYBZuAwVZFo5vT48+7PWYDTsBJfQ/QKqu/PcbDPndKt8zhnv8prrgA8JU
SOCN5DTY/CzFuE+/ajhCxJ035KeOcLlckwUHEixNIh0apV873YgHa31pIXNbOu8QVwNrNPIW5+ok
nqdN3bTIONHhYMu6/PeSdewRr3sN4zIeLOtnykJtecs0TNFFZLUwl7Q/NnAhjNlNv+ZLzs1RErjU
+1nVcopKtAD5HqD21v/HxWG/sMYkHo2EcHbXfYCbfUTJOasDm6qroh09ssbPE+LXZzCI3YfwWZlD
F23RcFtFD/yXS37OqVvWG1HwCnaxp+YwUqe76Z/JqUJrS8IoImKaWt0Zm+S5k/Yw3V+1qAjiKT7S
ODoFaf+hBWG2ZaZMT4FzO3jKx7zsA3reJYdrY3tk/n2PxPPX/U1dm1AEfKAZM6N64ZgMg+7eX4+w
8lwNCL9fr0ogrSLnlhqJzEB3wqjQYs+q4j+fB5/UNKW4VqSnTH8Tm1AWE7C25UnrP8ZOCBGzsoSD
h3/AK3NS7ru6nVaI9rHQRxms25lLx243TqEnZ0OBy+lELf1xBxmo35TU9g5fL0JESlHtRmFlBmnM
8mnFLx8R+T6H6p0sibXhRt6MsrFuX6UhLqCRCtqkEM8qjECqDZ4tzi1cpljM8JvqWw4qfe6NdNbi
UbxLYwLAN5CSxvt51T+54DgKvtTLZWOiwqUY3itStnRGJvumJp30K37Jy3TEbIXPOXLGyleyp9++
3Lh4F860xOcEWTJ4DQoGI0jKGYfMUpQ9IZJ89g+xvhPp+7iKfd33wsesydijNDNCLc/Q6Q6d3Y36
9X5bgmsJL3HnUGXQEXiHjIP9cUCrPcNCSYkJ4p615tIeKidB3pujtdJTE5pvqN2WbCqRTUTaH4+f
LFXvKkAEtVjho8qdMqIq6+E8OcRVYD2jWLoLA1BNthOcb6D0RojaBjH4YhFfK2LwRGBCTvWanxHt
akllA9HXXKLp+UjNI99cELTd07Cxdn9X8njd5YGKFX+g4FI2yzVBhLHE8vVuKpeyp0+Z/Rb+cwaL
QswlyDt6t56c80GUyG2r2wgcsKhJzlFWXqmbNvsz+DSN5j+gJZMmdVz6Ts/SJ+bpWigDrRlVmz8V
lV+InkOWn6LPywOvS/JiVEPaFEHOfUNxNk3+UKTCFF1DQFg+7Lb9qAsE5FKKXv2YvozA8UOeO0Gs
Fj7zTnFX241osNqBC1TWJcRlkUiRKqAJNf0+YcHYJGq05VSyXdfEVD8FRo0fFewLLmvepBydfahA
hvBrixGwELAr6Qti6NCDhN0Pj+2sRB6/YNon5UEUEgy6jTdD0lxHkvQsTHnh9HNU2I+ckVTG7b2Y
LHonCuO5GjGf9QyO6LTv+yR1ZqKPR2KWH7yFONynRD9jphgZDLYCFqzknSUoSYzMB7D+3U3GOWXK
b3Hh/N2Q39weDS0yzSDoICf44792/7zQaKDWAb7mf2oPQvatzmOpOeqg0oeKQzA9Gohvv4D8iPvc
kRlIjE4il2bCgHvaeXLowbBbj5+h1Mll2hXu/N5lgsuKW5D+Auh524+x/dwKDM6bgJrMZbB4Tezr
gGh0wbWF/Ao7zRVz2YmDPmTkAVZZV1WYaVfzpcL+PiAToIakhc/EiNlI+FxQRwguDzaBRv33vVWX
3gCFbU+pSg+lCeTAKpm5gVqClu+wJhVm4/7t+LJrHnnrQlegUSEj6Ccx2Pt5QcrkbG/QMW4=
`protect end_protected
